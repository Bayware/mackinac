package special_packet_pkg ;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "special_packet.svh"

endpackage 
