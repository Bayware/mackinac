// ===========================================================================================
// ===========================================================================================
// $File: 
//
// DESCRIPTION : 
// ===========================================================================================

`ifndef DEFINES 
`define DEFINES

`timescale 10ps/10ps

`define FLOW_LABEL_NBITS 20
`define IP_DA_NBITS 128
`define IP_SA_NBITS 128
`define VLAN_NBITS 16
`define MAC_NBITS 48

`define PACKET_LENGTH_NBITS             14
`define PACKET_LENGTH_RANGE             `PACKET_LENGTH_NBITS-1:0

`define RESET_SIG_DUP reset_dup_n
`define RESET_SIG reset_n
`define RESET_SIG_D1 reset_n_d1
`define ACTIVE_RESET ~reset_n
`define ACTIVE_RESET_LEVEL 1'b0
`define INACTIVE_RESET reset_n
`define INACTIVE_RESET_LEVEL 1'b1
`define COMBINE_RESET(R) ~(`ACTIVE_RESET|R)
`define RESET_EDGE negedge reset_n

`define RESET_SIG_AXI reset_axi_n
`define RESET_SIG_AXI_D1 reset_axi_n_d1
`define ACTIVE_RESET_AXI ~reset_axi_n
`define INACTIVE_RESET_AXI reset_axi_n
`define RESET_EDGE_AXI negedge reset_axi_n

`define RESET_SIG_MAC reset_mac_n
`define RESET_SIG_MAC_D1 reset_mac_n_d1
`define ACTIVE_RESET_MAC ~reset_mac_n
`define INACTIVE_RESET_MAC reset_mac_n
`define RESET_EDGE_MAC negedge reset_mac_n

`define SYNC_RST

`ifdef SYNC_RST
   `define CLK_RST posedge clk
   `define CLK_RST_AXI posedge clk_axi
   `define CLK_RST_MAC posedge clk_mac
`else 
   `define CLK_RST posedge clk or `RESET_EDGE
   `define CLK_RST_AXI posedge clk_axi or `RESET_EDGE_AXI
   `define CLK_RST_MAC posedge clk_mac or `RESET_EDGE_MAC
`endif

`define TIME_BASE_NBITS 10
`define REAL_TIME_NBITS 32

`define SUB_EXP_TIME_NBITS 16
`define EXP_TIME_NBITS 16

`define AGING_TIME_NBITS 10

`define DMA_BUS_NBITS          64

`define PORT_BUS_NBYTES          4
`define PORT_BUS_NBITS          32
`define PORT_BUS_RANGE          `PORT_BUS_NBITS-1:0
`define PORT_BUS_VB_NBITS          2
`define PORT_BUS_VB_RANGE          `PORT_BUS_VB_NBITS-1:0

`define DATA_PATH_NBYTES          16
`define DATA_PATH_NBITS          8*`DATA_PATH_NBYTES  
`define DATA_PATH_NBITS_PORT     8*4
`define DATA_PATH_RANGE          `DATA_PATH_NBITS-1:0  
`define DATA_PATH_VB_NBITS          4
`define DATA_PATH_VB_RANGE          `DATA_PATH_VB_NBITS-1:0

`define DATA_PATH_PORT_BUS_RATIO          `DATA_PATH_NBYTES/`PORT_BUS_NBYTES

`define EM_BUF_PTR_NBITS 12
`define EM_BUF_PTR_LSB_NBITS 2

`define BUF_SIZE             64 
`define BUF_SIZE_OVER_DATA_PATH_NBYTES             `BUF_SIZE/`DATA_PATH_NBYTES 

`define BUF_PTR_NBITS             12 
`define BUF_PTR_RANGE             `BUF_PTR_NBITS-1:0 
`define BUF_PTR_LSB_NBITS             2 
`define BUF_PTR_LSB_RANGE             `BUF_PTR_LSB_NBITS-1:0

`define PORT_ID_NBITS 3	
`define PORT_ID_RANGE `PORT_ID_NBITS-1:0	
`define NUM_OF_10G_PORTS 2   
`define NUM_OF_DMA_PORTS 4	
`define NUM_OF_OAM_PORTS 1	

`define NUM_OF_PORTS `NUM_OF_10G_PORTS+`NUM_OF_DMA_PORTS+`NUM_OF_OAM_PORTS

`define NUM_OF_PU 20
`define PU_ID_NBITS 5

`define NUM_OF_PIO 10

`define PIO_NBITS             32
`define PIO_ADDR_MSB             `PIO_NBITS-1
`define PIO_ADDR_LSB             0
`define PIO_ADDR_RANGE             `PIO_ADDR_MSB:`PIO_ADDR_LSB
`define PIO_RANGE             `PIO_NBITS-1:0


`define DISCARD_INFO_SRC_PORT_NBITS `PORT_ID_NBITS
`define DISCARD_INFO_LEN_NBITS `PACKET_LENGTH_NBITS
`define DISCARD_INFO_BUF_PTR_NBITS `BUF_PTR_NBITS
`define DISCARD_INFO_NBITS `DISCARD_INFO_SRC_PORT_NBITS+`DISCARD_INFO_LEN_NBITS+`DISCARD_INFO_BUF_PTR_NBITS
`define DISCARD_INFO_RANGE `DISCARD_INFO_NBITS-1:0
`define DISCARD_INFO_SRC_PORT_RANGE `DISCARD_INFO_SRC_PORT_NBITS-1:0
`define DISCARD_INFO_SRC_PORT_POS `DISCARD_INFO_SRC_PORT_NBITS-1
`define DISCARD_INFO_SRC_PORT `DISCARD_INFO_SRC_PORT_POS:0
`define DISCARD_INFO_LEN_RANGE `DISCARD_INFO_LEN_NBITS-1:0
`define DISCARD_INFO_LEN_POS `DISCARD_INFO_LEN_NBITS+`DISCARD_INFO_SRC_PORT_POS
`define DISCARD_INFO_LEN `DISCARD_INFO_LEN_POS:`DISCARD_INFO_SRC_PORT_POS+1
`define DISCARD_INFO_BUF_PTR_RANGE `DISCARD_INFO_BUF_PTR_NBITS-1:0
`define DISCARD_INFO_BUF_PTR_POS `DISCARD_INFO_BUF_PTR_NBITS+`DISCARD_INFO_LEN_POS
`define DISCARD_INFO_BUF_PTR `DISCARD_INFO_BUF_PTR_POS:`DISCARD_INFO_LEN_POS+1

`define PU_SWITCH_INFO 2'd0
`define PU_CONNECTION_CONTEXT 2'd1
`define PU_TAG_HASH_TABLE 2'd2
`define PU_TAG_VALUE 2'd3

`define SWITCH_INFO_DEPTH_NBITS 4
`define CONNECTION_CONTEXT_DEPTH_NBITS 6
`define TAG_RESULT_DEPTH_NBITS 3

`define PU_WIDTH_NBITS 32

`define PU_MEM_DEPTH_NBITS 32
`define PU_MEM_DEPTH_RANGE `PU_MEM_DEPTH_NBITS-1:1
`define PU_MEM_ADDRESSABLE_DEPTH_NBITS 20
`define PU_MEM_DEPTH_MSB_RANGE `PU_MEM_ADDRESSABLE_DEPTH_NBITS-1:`PU_MEM_ADDRESSABLE_DEPTH_NBITS-1-3
`define PU_MEM_DEPTH_LSB_RANGE `PU_MEM_DEPTH_NBITS-1-4:2
`define PU_PD_MEM 4'b0000
`define PU_RAS_MEM 4'b0001
`define PU_FLOW_MEM 4'b1000
`define PU_TOPIC_MEM 4'b1001
`define PU_SWITCH_INFO_MEM 4'b1010
`define PU_CONNECTION_CONTEXT_MEM 4'b1011
`define PU_TAG_LOOKUP_REQ 4'b1100
`define PU_TAG_LOOKUP_RESULT 4'b1101

`define PU_RAS_MEM_RAS 1'b0
`define PU_RAS_MEM_META 1'b1

`define PPL_LOC 0
`define PPL_NBITS 6
`define PPL_RANGE `PPL_NBITS-1:0
`define PPL_POS `DATA_PATH_NBITS-1-5*8-2
`define PPL `PPL_POS:`PPL_POS-`PPL_NBITS+1
`define ISSUER_ID_LOC 0
`define ISSUER_ID_NBITS 16
`define ISSUER_ID_RANGE `ISSUER_ID_NBITS-1:0
`define ISSUER_ID_POS `DATA_PATH_NBITS-1-6*8
`define ISSUER_ID `ISSUER_ID_POS:`ISSUER_ID_POS-`ISSUER_ID_NBITS+1
`define SERIAL_NUM_LOC 0
`define SERIAL_NUM_NBITS 64
`define SERIAL_NUM_RANGE `SERIAL_NUM_NBITS-1:0
`define SERIAL_NUM_POS `DATA_PATH_NBITS-1-8*8
`define SERIAL_NUM `SERIAL_NUM_POS:`SERIAL_NUM_POS-`SERIAL_NUM_NBITS+1
`define NOTAFTER_LOC 1
`define NOTAFTER_NBITS 16
`define NOTAFTER_RANGE `NOTAFTER_NBITS-1:0
`define NOTAFTER_POS `DATA_PATH_NBITS-1-4*8
`define NOTAFTER `NOTAFTER_POS:`NOTAFTER_POS-`NOTAFTER_NBITS+1
`define DOMAIN_ID_LOC 1
`define DOMAIN_ID_NBITS 24
`define DOMAIN_ID_RANGE `DOMAIN_ID_NBITS-1:0
`define DOMAIN_ID_POS `DATA_PATH_NBITS-1-8*8
`define DOMAIN_ID `DOMAIN_ID_POS:`DOMAIN_ID_POS-`DOMAIN_ID_NBITS+1
`define TOPIC_ROLE_LOC 1
`define TOPIC_ROLE_NBITS 8
`define TOPIC_ROLE_RANGE `TOPIC_ROLE_NBITS-1:0
`define TOPIC_ROLE_POS `DATA_PATH_NBITS-1-11*8
`define TOPIC_ROLE `TOPIC_ROLE_POS:`TOPIC_ROLE_POS-`TOPIC_ROLE_NBITS+1
`define MASKON_LOC 1
`define MASKON_NBITS 16
`define MASKON_RANGE `MASKON_NBITS-1:0
`define MASKON_POS `DATA_PATH_NBITS-1-12*8
`define MASKON `MASKON_POS:`MASKON_POS-`MASKON_NBITS+1
`define BA_LOC 1
`define BA_NBITS 6
`define BA_RANGE `BA_NBITS-1:0
`define BA_POS `DATA_PATH_NBITS-1-14*8
`define BA `BA_POS:`BA_POS-`BA_NBITS+1
`define EA_LOC 1
`define EA_NBITS 4
`define EA_RANGE `EA_NBITS-1:0
`define EA_POS `DATA_PATH_NBITS-1-14*8-`BA_NBITS
`define EA `EA_POS:`EA_POS-`EA_NBITS+1
`define FSPDA_LOC 1
`define FSPDA_NBITS 3
`define FSPDA_RANGE `FSPDA_NBITS-1:0
`define FSPDA_POS `DATA_PATH_NBITS-1-14*8-`BA_NBITS-`EA_NBITS
`define FSPDA `FSPDA_POS:`FSPDA_POS-`FSPDA_NBITS+1
`define TSPDA_LOC 1
`define TSPDA_NBITS 3
`define TSPDA_RANGE `TSPDA_NBITS-1:0
`define TSPDA_POS `DATA_PATH_NBITS-1-14*8-`BA_NBITS-`EA_NBITS-`FSPDA_NBITS
`define TSPDA `TSPDA_POS:`TSPDA_POS-`TSPDA_NBITS+1
`define SIGNATURE_LOC 2
`define SIGNATURE_NBITS 512
`define SIGNATURE_RANGE `SIGNATURE_NBITS-1:0
`define SIGNATURE_POS `DATA_PATH_NBITS-1

`define ECDSA_FLOW_ISSUER_ID_NBITS `ISSUER_ID_NBITS

`define STEP5D_FLOW_SERIAL_NUM_NBITS `SERIAL_NUM_NBITS

`define LOGIC_HASH_NBITS 256
`define TOPIC_POLICY_ROLE_NBITS (8+16)
`define TOPIC_POLICY_NBITS `TOPIC_POLICY_ROLE_NBITS*4

`define FLOW_LH_PPL_NBITS `PPL_NBITS

`define FLOW_PU_MASKON_NBITS 2
`define FLOW_PU_EA_NBITS `EA_NBITS
`define FLOW_PU_FSPDA_NBITS `FSPDA_NBITS
`define FLOW_PU_TSPDA_NBITS `TSPDA_NBITS
`define FLOW_PU_NBITS `FLOW_PU_MASKON_NBITS+`FLOW_PU_EA_NBITS+`FLOW_PU_FSPDA_NBITS+`FLOW_PU_TSPDA_NBITS
`define FLOW_PU_RANGE `FLOW_PU_NBITS-1:0
`define FLOW_PU_MASKON_RANGE `FLOW_PU_MASKON_NBITS-1:0
`define FLOW_PU_MASKON_POS `FLOW_PU_MASKON_NBITS-1
`define FLOW_PU_MASKON `FLOW_PU_MASKON_POS:0
`define FLOW_PU_EA_RANGE `FLOW_PU_EA_NBITS-1:0
`define FLOW_PU_EA_POS `FLOW_PU_EA_NBITS+`FLOW_PU_MASKON_POS
`define FLOW_PU_EA `FLOW_PU_EA_POS:`FLOW_PU_MASKON_POS+1
`define FLOW_PU_FSPDA_RANGE `FLOW_PU_FSPDA_NBITS-1:0
`define FLOW_PU_FSPDA_POS `FLOW_PU_FSPDA_NBITS+`FLOW_PU_EA_POS
`define FLOW_PU_FSPDA `FLOW_PU_FSPDA_POS:`FLOW_PU_EA_POS+1
`define FLOW_PU_TSPDA_RANGE `FLOW_PU_TSPDA_NBITS-1:0
`define FLOW_PU_TSPDA_POS `FLOW_PU_TSPDA_NBITS+`FLOW_PU_FSPDA_POS
`define FLOW_PU_TSPDA `FLOW_PU_TSPDA_POS:`FLOW_PU_FSPDA_POS+1

`define FLOW_VALUE_IP_DA_NBITS `IP_DA_NBITS
`define FLOW_VALUE_IP_SA_NBITS `IP_SA_NBITS
`define FLOW_VALUE_FLOW_LABEL_NBITS `FLOW_LABEL_NBITS
`define FLOW_VALUE_NBITS `FLOW_VALUE_FLOW_LABEL_NBITS+`FLOW_VALUE_IP_SA_NBITS+`FLOW_VALUE_IP_DA_NBITS
`define FLOW_VALUE_RANGE `FLOW_VALUE_NBITS-1:0
`define FLOW_VALUE_IP_DA_RANGE `FLOW_VALUE_IP_DA_NBITS-1:0
`define FLOW_VALUE_IP_DA_POS `FLOW_VALUE_IP_DA_NBITS-1
`define FLOW_VALUE_IP_DA `FLOW_VALUE_IP_DA_POS:0
`define FLOW_VALUE_IP_SA_RANGE `FLOW_VALUE_IP_SA_NBITS-1:0
`define FLOW_VALUE_IP_SA_POS `FLOW_VALUE_IP_SA_NBITS+`FLOW_VALUE_IP_DA_POS
`define FLOW_VALUE_IP_SA `FLOW_VALUE_IP_SA_POS:`FLOW_VALUE_IP_DA_POS+1
`define FLOW_VALUE_FLOW_LABEL_RANGE `FLOW_VALUE_FLOW_LABEL_NBITS-1:0
`define FLOW_VALUE_FLOW_LABEL_POS `FLOW_VALUE_FLOW_LABEL_NBITS+`FLOW_VALUE_IP_SA_POS
`define FLOW_VALUE_FLOW_LABEL `FLOW_VALUE_FLOW_LABEL_POS:`FLOW_VALUE_IP_SA_POS+1

`define FLOW_NUM_OF_ENTRIES 2
`define FLOW_NUM_OF_ENTRIES_NBITS 1
`define FLOW_NUM_OF_HASH TABLES 2
`define FLOW_NUM_OF_HASH_TABLES_NBITS 1

`define FID_NBITS 12
`define FID_RANGE `FID_NBITS-1:0
`define TID_NBITS 10

`define FLOW_KEY_NBITS (`IP_SA_NBITS+`IP_DA_NBITS+`FLOW_LABEL_NBITS)
`define FLOW_VALUE_DEPTH_NBITS `FID_NBITS
`define FLOW_HASH_TABLE_DEPTH_NBITS (`FLOW_VALUE_DEPTH_NBITS-`FLOW_NUM_OF_HASH_TABLES_NBITS-`FLOW_NUM_OF_ENTRIES_NBITS)
`define FLOW_HASH_ENTRY_NBITS (`FLOW_VALUE_DEPTH_NBITS+`FLOW_HASH_TABLE_DEPTH_NBITS)
`define FLOW_HASH_BUCKET_NBITS `FLOW_HASH_ENTRY_NBITS*`FLOW_NUM_OF_ENTRIES
`define FLOW_VALUE_KEY `FLOW_KEY_NBITS-1:0

`define SWITCH_TAG_NBITS 8

`define TOPIC_NUM_OF_ENTRIES 2
`define TOPIC_NUM_OF_ENTRIES_NBITS 1
`define TOPIC_NUM_OF_HASH TABLES 2
`define TOPIC_NUM_OF_HASH_TABLES_NBITS 1

`define TOPIC_KEY_NBITS `IP_DA_NBITS
`define TOPIC_VALUE_DEPTH_NBITS `TID_NBITS
`define TOPIC_HASH_TABLE_DEPTH_NBITS (`TOPIC_VALUE_DEPTH_NBITS-`TOPIC_NUM_OF_HASH_TABLES_NBITS-`TOPIC_NUM_OF_ENTRIES_NBITS)
`define TOPIC_HASH_ENTRY_NBITS (`TOPIC_VALUE_DEPTH_NBITS+`TOPIC_HASH_TABLE_DEPTH_NBITS)
`define TOPIC_HASH_BUCKET_NBITS (`TOPIC_HASH_ENTRY_NBITS*`TOPIC_NUM_OF_ENTRIES)
`define TOPIC_VALUE_KEY `TOPIC_KEY_NBITS-1:0
`define TOPIC_VALUE_NBITS `TOPIC_KEY_NBITS

`define ASA_RCI2SCI_TABLE             6'd0

`define ENCRYPTION_KEY_NBITS 256

`define SPI_NBITS 32
`define SEQUENCE_NUMBER_NBITS 32

`define TRAFFIC_CLASS_NBITS 8	
`define PRI_NBITS 3	
`define RCI_NBITS 13
`define RCI_TYPE_NBITS 3
`define HOP_NBITS `RCI_NBITS+`RCI_TYPE_NBITS
`define SCI_NBITS 6	
`define PACKET_ID_NBITS `SCI_NBITS	
`define SCI_VEC_NBITS (1<<`SCI_NBITS)	
`define DEFAULT_RCI 16'h0a

`define EKEY_NUM_OF_ENTRIES 2
`define EKEY_NUM_OF_ENTRIES_NBITS 1
`define EKEY_NUM_OF_HASH TABLES 2
`define EKEY_NUM_OF_HASH_TABLES_NBITS 1

`define EKEY_KEY_NBITS `SPI_NBITS
`define EKEY_VALUE_DEPTH_NBITS 9
`define EKEY_VALUE_NBITS (`SEQUENCE_NUMBER_NBITS+`EKEY_KEY_NBITS+`ENCRYPTION_KEY_NBITS)
`define EKEY_HASH_TABLE_DEPTH_NBITS (`EKEY_VALUE_DEPTH_NBITS-`EKEY_NUM_OF_HASH_TABLES_NBITS-`EKEY_NUM_OF_ENTRIES_NBITS)
`define EKEY_HASH_ENTRY_NBITS (1+`EKEY_VALUE_DEPTH_NBITS+`EKEY_HASH_TABLE_DEPTH_NBITS)
`define EKEY_HASH_BUCKET_NBITS (`EKEY_HASH_ENTRY_NBITS*`EKEY_NUM_OF_ENTRIES)
`define EKEY_VALUE_KEY `EKEY_KEY_NBITS-1:0
`define EKEY_VALUE_SN `SEQUENCE_NUMBER_NBITS+`EKEY_KEY_NBITS-1:`EKEY_KEY_NBITS
`define EKEY_VALUE_PAYLOAD `EKEY_VALUE_NBITS-1:`SEQUENCE_NUMBER_NBITS+`EKEY_KEY_NBITS

`define RCI_NUM_OF_ENTRIES 2
`define RCI_NUM_OF_ENTRIES_NBITS 1
`define RCI_NUM_OF_HASH TABLES 2
`define RCI_NUM_OF_HASH_TABLES_NBITS 1

`define RCI_KEY_NBITS 256
`define RCI_VALUE_DEPTH_NBITS 6
`define RCI_VALUE_NBITS `RCI_KEY_NBITS+`RCI_NBITS
`define RCI_HASH_TABLE_DEPTH_NBITS (`RCI_VALUE_DEPTH_NBITS-`RCI_NUM_OF_HASH_TABLES_NBITS-`RCI_NUM_OF_ENTRIES_NBITS)
`define RCI_HASH_ENTRY_NBITS (1+`RCI_VALUE_DEPTH_NBITS+`RCI_HASH_TABLE_DEPTH_NBITS)
`define RCI_HASH_BUCKET_NBITS (`RCI_HASH_ENTRY_NBITS*`RCI_NUM_OF_ENTRIES)
`define RCI_VALUE_KEY `RCI_KEY_NBITS-1:0
`define RCI_VALUE_PAYLOAD `RCI_VALUE_NBITS-1:`RCI_KEY_NBITS

`define EEKEY_NUM_OF_ENTRIES 2
`define EEKEY_NUM_OF_ENTRIES_NBITS 1
`define EEKEY_NUM_OF_HASH TABLES 2
`define EEKEY_NUM_OF_HASH_TABLES_NBITS 1

`define EEKEY_KEY_NBITS `SPI_NBITS
`define EEKEY_VALUE_DEPTH_NBITS 9
`define EEKEY_VALUE_PAYLOAD_NBITS (`SEQUENCE_NUMBER_NBITS+`ENCRYPTION_KEY_NBITS)
`define EEKEY_VALUE_NBITS (`EEKEY_VALUE_PAYLOAD_NBITS+`EEKEY_KEY_NBITS)
`define EEKEY_HASH_TABLE_DEPTH_NBITS (`EEKEY_VALUE_DEPTH_NBITS-`EEKEY_NUM_OF_HASH_TABLES_NBITS-`EEKEY_NUM_OF_ENTRIES_NBITS)
`define EEKEY_HASH_ENTRY_NBITS (1+`EEKEY_VALUE_DEPTH_NBITS+`EEKEY_HASH_TABLE_DEPTH_NBITS)
`define EEKEY_HASH_BUCKET_NBITS (`EEKEY_HASH_ENTRY_NBITS*`EEKEY_NUM_OF_ENTRIES)
`define EEKEY_VALUE_KEY `EEKEY_KEY_NBITS-1:0
`define EEKEY_VALUE_SN `SEQUENCE_NUMBER_NBITS+`EEKEY_KEY_NBITS-1:`EEKEY_KEY_NBITS
`define EEKEY_VALUE_EKEY EEKEY_VALUE_NBITS-1:`SEQUENCE_NUMBER_NBITS+`EEKEY_KEY_NBITS
`define EEKEY_VALUE_PAYLOAD `EEKEY_VALUE_NBITS-1:`EEKEY_KEY_NBITS

`define TUNNEL_NUM_OF_ENTRIES 2
`define TUNNEL_NUM_OF_ENTRIES_NBITS 1
`define TUNNEL_NUM_OF_HASH TABLES 2
`define TUNNEL_NUM_OF_HASH_TABLES_NBITS 1

`define TUNNEL_KEY_NBITS `RCI_NBITS
`define TUNNEL_VALUE_DEPTH_NBITS 6
`define TUNNEL_HASH_TABLE_DEPTH_NBITS (`TUNNEL_VALUE_DEPTH_NBITS-`TUNNEL_NUM_OF_HASH_TABLES_NBITS-`TUNNEL_NUM_OF_ENTRIES_NBITS)
`define TUNNEL_HASH_ENTRY_NBITS (1+`TUNNEL_VALUE_DEPTH_NBITS+`TUNNEL_HASH_TABLE_DEPTH_NBITS)
`define TUNNEL_HASH_BUCKET_NBITS (`TUNNEL_HASH_ENTRY_NBITS*`TUNNEL_NUM_OF_ENTRIES)

`define TUNNEL_VALUE_KEY_NBITS `TUNNEL_KEY_NBITS
`define TUNNEL_VALUE_KEY_RANGE `TUNNEL_VALUE_KEY_NBITS-1:0
`define TUNNEL_VALUE_KEY_POS `TUNNEL_VALUE_KEY_NBITS-1
`define TUNNEL_VALUE_KEY `TUNNEL_VALUE_KEY_POS:0

`define TUNNEL_VALUE_IP_DA_NBITS `IP_DA_NBITS
`define TUNNEL_VALUE_IP_SA_NBITS `IP_SA_NBITS
`define TUNNEL_VALUE_VLAN_NBITS `VLAN_NBITS
`define TUNNEL_VALUE_MAC_NBITS `MAC_NBITS
`define TUNNEL_VALUE_SPI_NBITS `SPI_NBITS
`define TUNNEL_VALUE_SN_NBITS `SERIAL_NUM_NBITS
`define TUNNEL_VALUE_PAYLOAD_NBITS (`TUNNEL_VALUE_VLAN_NBITS+`TUNNEL_VALUE_IP_SA_NBITS+`TUNNEL_VALUE_IP_DA_NBITS+`TUNNEL_VALUE_MAC_NBITS+`TUNNEL_VALUE_SPI_NBITS+`TUNNEL_VALUE_SN_NBITS)
`define TUNNEL_VALUE_RANGE `TUNNEL_VALUE_NBITS-1:0
`define TUNNEL_VALUE_IP_DA_RANGE `TUNNEL_VALUE_IP_DA_NBITS-1:0
`define TUNNEL_VALUE_IP_DA_POS `TUNNEL_VALUE_IP_DA_NBITS-1
`define TUNNEL_VALUE_IP_DA `TUNNEL_VALUE_IP_DA_POS:0
`define TUNNEL_VALUE_IP_SA_RANGE `TUNNEL_VALUE_IP_SA_NBITS-1:0
`define TUNNEL_VALUE_IP_SA_POS `TUNNEL_VALUE_IP_SA_NBITS+`TUNNEL_VALUE_IP_DA_POS
`define TUNNEL_VALUE_IP_SA `TUNNEL_VALUE_IP_SA_POS:`TUNNEL_VALUE_IP_DA_POS+1
`define TUNNEL_VALUE_VLAN_RANGE `TUNNEL_VALUE_VLAN_NBITS-1:0
`define TUNNEL_VALUE_VLAN_POS `TUNNEL_VALUE_VLAN_NBITS+`TUNNEL_VALUE_IP_SA_POS
`define TUNNEL_VALUE_VLAN `TUNNEL_VALUE_VLAN_POS:`TUNNEL_VALUE_IP_SA_POS+1
`define TUNNEL_VALUE_MAC_RANGE `TUNNEL_VALUE_MAC_NBITS-1:0
`define TUNNEL_VALUE_MAC_POS `TUNNEL_VALUE_MAC_NBITS+`TUNNEL_VALUE_VLAN_POS
`define TUNNEL_VALUE_MAC `TUNNEL_VALUE_MAC_POS:`TUNNEL_VALUE_VLAN_POS+1
`define TUNNEL_VALUE_SPI_RANGE `TUNNEL_VALUE_SPI_NBITS-1:0
`define TUNNEL_VALUE_SPI_POS `TUNNEL_VALUE_SPI_NBITS+`TUNNEL_VALUE_MAC_POS
`define TUNNEL_VALUE_SPI `TUNNEL_VALUE_SPI_POS:`TUNNEL_VALUE_MAC_POS+1
`define TUNNEL_VALUE_SN_RANGE `TUNNEL_VALUE_SN_NBITS-1:0
`define TUNNEL_VALUE_SN_POS `TUNNEL_VALUE_SN_NBITS+`TUNNEL_VALUE_SPI_POS
`define TUNNEL_VALUE_SN `TUNNEL_VALUE_SN_POS:`TUNNEL_VALUE_SPI_POS+1

`define TUNNEL_VALUE_NBITS (`TUNNEL_VALUE_PAYLOAD_NBITS+`TUNNEL_VALUE_KEY_NBITS)
`define TUNNEL_VALUE_PAYLOAD `TUNNEL_VALUE_NBITS-1:`TUNNEL_VALUE_KEY_NBITS


`define TAG_NBITS 24

`define TAG_NUM_OF_ENTRIES 4
`define TAG_NUM_OF_ENTRIES_NBITS 2
`define TAG_NUM_OF_HASH TABLES 2
`define TAG_NUM_OF_HASH_TABLES_NBITS 1

`define TAG_KEY_NBITS `TAG_NBITS
`define TAG_VALUE_DEPTH_NBITS 8
`define TAG_HASH_TABLE_DEPTH_NBITS (`TAG_VALUE_DEPTH_NBITS-`TAG_NUM_OF_HASH_TABLES_NBITS-`TAG_NUM_OF_ENTRIES_NBITS)
`define TAG_HASH_ENTRY_NBITS (`TAG_VALUE_DEPTH_NBITS+`TAG_HASH_TABLE_DEPTH_NBITS)
`define TAG_HASH_BUCKET_NBITS (`TAG_HASH_ENTRY_NBITS*`TAG_NUM_OF_ENTRIES)

`define TAG_VALUE_PAYLOAD_NBITS `RCI_NBITS
`define TAG_VALUE_NBITS (`RCI_NBITS+`TAG_KEY_NBITS)
`define TAG_VALUE_PAYLOAD `TAG_VALUE_NBITS-1:`TAG_KEY_NBITS
`define TAG_VALUE_KEY `TAG_KEY_NBITS-1:0

`define PIARB_BUF_PTR_NBITS 12
`define PIARB_BUF_PTR_LSB_NBITS 1
`define PIARB_INST_BUF_PTR_NBITS 12
`define PIARB_INST_BUF_PTR_LSB_NBITS 1
`define PU_QUEUE_ENTRIES_NBITS 11

`define INITIAL_HOP 16'hFFFF

`define PP_PU_FIFO_DEPTH_NBITS 6	
`define HOP_INFO_FIFO_DEPTH_NBITS 6	

`define PROC_LEV_NBITS 6	
`define PROC_LEV_RANGE `PROC_LEV_NBITS-1:0	

`define HOP_DESC_NBITS 6	
`define HOP_ID_NBITS 6	
`define HOP_ID_RANGE `HOP_IP_NBITS-1:0	

`define PIARB_BUF_FIFO_DEPTH_NBITS 7
`define PIARB_INST_BUF_FIFO_DEPTH_NBITS 8

`define CHUNK_TYPE_NBITS 4
`define CHUNK_LEN_NBITS 12

`define PATH_CHUNK_NBITS 7
`define INST_CHUNK_NBITS 11
`define PD_CHUNK_NBITS 7

`define PATH_CHUNK_NBYTES        256
`define PATH_CHUNK_DEPTH        (`PATH_CHUNK_NBYTES/`DATA_PATH_NBYTES)
`define PATH_CHUNK_DEPTH_NBITS  4
`define PATH_CHUNK_ADDR_RANGE  `PATH_CHUNK_DEPTH_NBITS:0

`define PD_CHUNK_NBYTES        128
`define PD_CHUNK_DEPTH_NBITS  7

`define TOPIC_PD_NBITS 6
`define FLOW_PD_NBITS 6

`define SP_HEADER_LENGTH_UNIT       8
`define SP_HEADER_LENGTH_NBITS       8
`define HEADER_LENGTH        (((1<<SP_HEADER_LENGTH_NBITS)*`SP_HEADER_LENGTH_UNIT+48)/`DATA_PATH_NBYTES)
`define HEADER_LENGTH_NBITS  (`CHUNK_LEN_NBITS+2-4)
`define HEADER_LENGTH_RANGE  `HEADER_LENGTH_NBITS-1:0

`define CIR_NBITS 16
`define EIR_NBITS 16

`define LIMITER_NBITS `BA_NBITS
`define LIMITING_PROFILE_NBITS (`CIR_NBITS<<1)

`define FILL_TB_NBITS (`PORT_ID_NBITS+`LIMITER_NBITS)

`define TQNA_NBITS 16
`define WDRR_QUANTUM_NBITS 16
`define WDRR_N_NBITS 16
`define SHAPING_PROFILE_NBITS (`CIR_NBITS<<1)
`define DEFICIT_COUNTER_NBITS 16

`define FIRST_LVL_SCH_ID_NBITS 7
`define SECOND_LVL_SCH_ID_NBITS 5
`define THIRD_LVL_SCH_ID_NBITS 4
`define FOURTH_LVL_SCH_ID_NBITS 3	
	
// 1st: 256; 2nd: 128; 3rd: 28, 4th: 14
`define FIRST_LVL_QUEUE_ID_NBITS	8
`define SECOND_LVL_QUEUE_ID_NBITS `FIRST_LVL_SCH_ID_NBITS
`define THIRD_LVL_QUEUE_ID_NBITS `SECOND_LVL_SCH_ID_NBITS
`define FOURTH_LVL_QUEUE_ID_NBITS `THIRD_LVL_SCH_ID_NBITS

`define FIRST_LVL_QUEUE_PROFILE_NBITS	(4+`FIRST_LVL_SCH_ID_NBITS)
`define SECOND_LVL_QUEUE_PROFILE_NBITS	(4+`SECOND_LVL_SCH_ID_NBITS)
`define THIRD_LVL_QUEUE_PROFILE_NBITS	(4+`THIRD_LVL_SCH_ID_NBITS)
`define FOURTH_LVL_QUEUE_PROFILE_NBITS	(4+`FOURTH_LVL_SCH_ID_NBITS)

`define QUEUE_ASSOCIATION_NBITS (`PORT_ID_NBITS+`FOURTH_LVL_QUEUE_ID_NBITS+`THIRD_LVL_QUEUE_ID_NBITS+`SECOND_LVL_QUEUE_ID_NBITS)

`define READ_COUNT_NBITS 6	
`define READ_COUNT_RANGE `READ_COUNT_NBITS-1:0	

`define PU_ASA_TS_NBITS 3
`define PU_ASA_TS 7
`define PU_ASA_NBITS 32

`define ACTION_SET_TYPE_NBITS 2

`define FLOW_ACTION_NBITS (`SCI_VEC_NBITS+`ACTION_SET_TYPE_NBITS)

`define FLOW_POLICY2_TCLASS_NBITS `TRAFFIC_CLASS_NBITS
`define FLOW_POLICY2_DOMAIN_ID_NBITS `DOMAIN_ID_NBITS
`define FLOW_POLICY2_MASKON_NBITS `MASKON_NBITS-6
`define FLOW_POLICY2_NBITS (`FLOW_POLICY2_MASKON_NBITS+`FLOW_POLICY2_DOMAIN_ID_NBITS+`FLOW_POLICY2_TCLASS_NBITS)
`define FLOW_POLICY2_RANGE `FLOW_POLICY2_NBITS-1:0
`define FLOW_POLICY2_TCLASS_RANGE `FLOW_POLICY2_TCLASS_NBITS-1:0
`define FLOW_POLICY2_TCLASS_POS `FLOW_POLICY2_TCLASS_NBITS-1
`define FLOW_POLICY2_TCLASS `FLOW_POLICY2_TCLASS_POS:0
`define FLOW_POLICY2_DOMAIN_ID_RANGE `FLOW_POLICY2_DOMAIN_ID_NBITS-1:0
`define FLOW_POLICY2_DOMAIN_ID_POS (`FLOW_POLICY2_DOMAIN_ID_NBITS+`FLOW_POLICY2_TCLASS_POS)
`define FLOW_POLICY2_DOMAIN_ID `FLOW_POLICY2_DOMAIN_ID_POS:`FLOW_POLICY2_TCLASS_POS+1
`define FLOW_POLICY2_MASKON_RANGE `FLOW_POLICY2_MASKON_NBITS-1:0
`define FLOW_POLICY2_MASKON_POS (`FLOW_POLICY2_MASKON_NBITS+`FLOW_POLICY2_DOMAIN_ID_POS)
`define FLOW_POLICY2_MASKON `FLOW_POLICY2_MASKON_POS:`FLOW_POLICY2_DOMAIN_ID_POS+1

`define AGGR_PAR_META_HDR_LEN_NBITS `HEADER_LENGTH_NBITS
`define AGGR_PAR_META_BUF_PTR_NBITS `BUF_PTR_NBITS
`define AGGR_PAR_META_LEN_NBITS `PACKET_LENGTH_NBITS
`define AGGR_PAR_META_PORT_NBITS `PORT_ID_NBITS
`define AGGR_PAR_META_RCI_NBITS `RCI_NBITS
`define AGGR_PAR_META_DISCARD_NBITS 1
`define AGGR_PAR_META_NBITS (`AGGR_PAR_META_LEN_NBITS+`AGGR_PAR_META_BUF_PTR_NBITS+`AGGR_PAR_META_HDR_LEN_NBITS+`AGGR_PAR_META_PORT_NBITS+`AGGR_PAR_META_RCI_NBITS+`AGGR_PAR_META_DISCARD_NBITS)
`define AGGR_PAR_META_RANGE `AGGR_PAR_META_NBITS-1:0
`define AGGR_PAR_META_HDR_LEN_RANGE `AGGR_PAR_META_HDR_LEN_NBITS-1:0
`define AGGR_PAR_META_HDR_LEN_POS `AGGR_PAR_META_HDR_LEN_NBITS-1
`define AGGR_PAR_META_HDR_LEN `AGGR_PAR_META_HDR_LEN_POS:0
`define AGGR_PAR_META_BUF_PTR_RANGE `AGGR_PAR_META_BUF_PTR_NBITS-1:0
`define AGGR_PAR_META_BUF_PTR_POS (`AGGR_PAR_META_BUF_PTR_NBITS+`AGGR_PAR_META_HDR_LEN_POS)
`define AGGR_PAR_META_BUF_PTR `AGGR_PAR_META_BUF_PTR_POS:`AGGR_PAR_META_HDR_LEN_POS+1
`define AGGR_PAR_META_LEN_RANGE `AGGR_PAR_META_LEN_NBITS-1:0
`define AGGR_PAR_META_LEN_POS `AGGR_PAR_META_LEN_NBITS+`AGGR_PAR_META_BUF_PTR_POS
`define AGGR_PAR_META_LEN `AGGR_PAR_META_LEN_POS:`AGGR_PAR_META_BUF_PTR_POS+1
`define AGGR_PAR_META_PORT_RANGE `AGGR_PAR_META_PORT_NBITS-1:0
`define AGGR_PAR_META_PORT_POS `AGGR_PAR_META_PORT_NBITS+`AGGR_PAR_META_LEN_POS
`define AGGR_PAR_META_PORT `AGGR_PAR_META_PORT_POS:`AGGR_PAR_META_LEN_POS+1
`define AGGR_PAR_META_RCI_RANGE `AGGR_PAR_META_RCI_NBITS-1:0
`define AGGR_PAR_META_RCI_POS `AGGR_PAR_META_RCI_NBITS+`AGGR_PAR_META_PORT_POS
`define AGGR_PAR_META_RCI `AGGR_PAR_META_RCI_POS:`AGGR_PAR_META_PORT_POS+1
`define AGGR_PAR_META_DISCARD_RANGE `AGGR_PAR_META_DISCARD_NBITS-1:0
`define AGGR_PAR_META_DISCARD_POS `AGGR_PAR_META_DISCARD_NBITS+`AGGR_PAR_META_RCI_POS
`define AGGR_PAR_META_DISCARD `AGGR_PAR_META_DISCARD_POS:`AGGR_PAR_META_RCI_POS+1

`define CLA_IRL_META_TRAFFIC_CLASS_NBITS `TRAFFIC_CLASS_NBITS
`define CLA_IRL_META_HDR_LEN_NBITS `HEADER_LENGTH_NBITS
`define CLA_IRL_META_BUF_PTR_NBITS `BUF_PTR_NBITS
`define CLA_IRL_META_LEN_NBITS `PACKET_LENGTH_NBITS
`define CLA_IRL_META_PORT_NBITS `PORT_ID_NBITS
`define CLA_IRL_META_RCI_NBITS `RCI_NBITS
`define CLA_IRL_META_FID_NBITS `FID_NBITS
`define CLA_IRL_META_TID_NBITS `TID_NBITS
`define CLA_IRL_META_TYPE1_NBITS 1
`define CLA_IRL_META_TYPE3_NBITS 1
`define CLA_IRL_META_DISCARD_NBITS 1
`define CLA_IRL_META_NBITS `CLA_IRL_META_TRAFFIC_CLASS_NBITS+`CLA_IRL_META_LEN_NBITS+`CLA_IRL_META_BUF_PTR_NBITS+`CLA_IRL_META_HDR_LEN_NBITS+`CLA_IRL_META_PORT_NBITS+`CLA_IRL_META_RCI_NBITS+`CLA_IRL_META_FID_NBITS+`CLA_IRL_META_TID_NBITS+`CLA_IRL_META_TYPE1_NBITS+`CLA_IRL_META_TYPE3_NBITS+`CLA_IRL_META_DISCARD_NBITS
`define CLA_IRL_META_RANGE `CLA_IRL_META_NBITS-1:0
`define CLA_IRL_META_TRAFFIC_CLASS_RANGE `CLA_IRL_META_TRAFFIC_CLASS_NBITS-1:0
`define CLA_IRL_META_TRAFFIC_CLASS_POS `CLA_IRL_META_TRAFFIC_CLASS_NBITS-1
`define CLA_IRL_META_TRAFFIC_CLASS `CLA_IRL_META_TRAFFIC_CLASS_POS:0
`define CLA_IRL_META_HDR_LEN_RANGE `CLA_IRL_META_HDR_LEN_NBITS-1:0
`define CLA_IRL_META_HDR_LEN_POS `CLA_IRL_META_HDR_LEN_NBITS+`CLA_IRL_META_TRAFFIC_CLASS_POS
`define CLA_IRL_META_HDR_LEN `CLA_IRL_META_HDR_LEN_POS:`CLA_IRL_META_TRAFFIC_CLASS_POS+1
`define CLA_IRL_META_BUF_PTR_RANGE `CLA_IRL_META_BUF_PTR_NBITS-1:0
`define CLA_IRL_META_BUF_PTR_POS `CLA_IRL_META_BUF_PTR_NBITS+`CLA_IRL_META_HDR_LEN_POS
`define CLA_IRL_META_BUF_PTR `CLA_IRL_META_BUF_PTR_POS:`CLA_IRL_META_HDR_LEN_POS+1
`define CLA_IRL_META_LEN_RANGE `CLA_IRL_META_LEN_NBITS-1:0
`define CLA_IRL_META_LEN_POS `CLA_IRL_META_LEN_NBITS+`CLA_IRL_META_BUF_PTR_POS
`define CLA_IRL_META_LEN `CLA_IRL_META_LEN_POS:`CLA_IRL_META_BUF_PTR_POS+1
`define CLA_IRL_META_PORT_RANGE `CLA_IRL_META_PORT_NBITS-1:0
`define CLA_IRL_META_PORT_POS `CLA_IRL_META_PORT_NBITS+`CLA_IRL_META_LEN_POS
`define CLA_IRL_META_PORT `CLA_IRL_META_PORT_POS:`CLA_IRL_META_LEN_POS+1
`define CLA_IRL_META_RCI_RANGE `CLA_IRL_META_RCI_NBITS-1:0
`define CLA_IRL_META_RCI_POS `CLA_IRL_META_RCI_NBITS+`CLA_IRL_META_PORT_POS
`define CLA_IRL_META_RCI `CLA_IRL_META_RCI_POS:`CLA_IRL_META_PORT_POS+1
`define CLA_IRL_META_FID_RANGE `CLA_IRL_META_FID_NBITS-1:0
`define CLA_IRL_META_FID_POS `CLA_IRL_META_FID_NBITS+`CLA_IRL_META_RCI_POS
`define CLA_IRL_META_FID `CLA_IRL_META_FID_POS:`CLA_IRL_META_RCI_POS+1
`define CLA_IRL_META_TID_RANGE `CLA_IRL_META_TID_NBITS-1:0
`define CLA_IRL_META_TID_POS `CLA_IRL_META_TID_NBITS+`CLA_IRL_META_FID_POS
`define CLA_IRL_META_TID `CLA_IRL_META_TID_POS:`CLA_IRL_META_FID_POS+1
`define CLA_IRL_META_TYPE1_RANGE `CLA_IRL_META_TYPE1_NBITS-1:0
`define CLA_IRL_META_TYPE1_POS `CLA_IRL_META_TYPE1_NBITS+`CLA_IRL_META_TID_POS
`define CLA_IRL_META_TYPE1 `CLA_IRL_META_TYPE1_POS:`CLA_IRL_META_TID_POS+1
`define CLA_IRL_META_TYPE3_RANGE `CLA_IRL_META_TYPE3_NBITS-1:0
`define CLA_IRL_META_TYPE3_POS `CLA_IRL_META_TYPE3_NBITS+`CLA_IRL_META_TYPE1_POS
`define CLA_IRL_META_TYPE3 `CLA_IRL_META_TYPE3_POS:`CLA_IRL_META_TYPE1_POS+1
`define CLA_IRL_META_DISCARD_RANGE `CLA_IRL_META_DISCARD_NBITS-1:0
`define CLA_IRL_META_DISCARD_POS `CLA_IRL_META_DISCARD_NBITS+`CLA_IRL_META_TYPE3_POS
`define CLA_IRL_META_DISCARD `CLA_IRL_META_DISCARD_POS:`CLA_IRL_META_TYPE3_POS+1

`define IRL_LH_META_TRAFFIC_CLASS_NBITS `TRAFFIC_CLASS_NBITS
`define IRL_LH_META_HDR_LEN_NBITS `HEADER_LENGTH_NBITS
`define IRL_LH_META_BUF_PTR_NBITS `BUF_PTR_NBITS
`define IRL_LH_META_LEN_NBITS `PACKET_LENGTH_NBITS
`define IRL_LH_META_PORT_NBITS `PORT_ID_NBITS
`define IRL_LH_META_RCI_NBITS `RCI_NBITS
`define IRL_LH_META_FID_NBITS `FID_NBITS
`define IRL_LH_META_TID_NBITS `TID_NBITS
`define IRL_LH_META_TYPE1_NBITS 1
`define IRL_LH_META_TYPE3_NBITS 1
`define IRL_LH_META_DISCARD_NBITS 1
`define IRL_LH_META_NBITS `IRL_LH_META_TRAFFIC_CLASS_NBITS+`IRL_LH_META_LEN_NBITS+`IRL_LH_META_BUF_PTR_NBITS+`IRL_LH_META_HDR_LEN_NBITS+`IRL_LH_META_PORT_NBITS+`IRL_LH_META_RCI_NBITS+`IRL_LH_META_FID_NBITS+`IRL_LH_META_TID_NBITS+`IRL_LH_META_TYPE1_NBITS+`IRL_LH_META_TYPE3_NBITS+`IRL_LH_META_DISCARD_NBITS
`define IRL_LH_META_RANGE `IRL_LH_META_NBITS-1:0
`define IRL_LH_META_TRAFFIC_CLASS_RANGE `IRL_LH_META_TRAFFIC_CLASS_NBITS-1:0
`define IRL_LH_META_TRAFFIC_CLASS_POS `IRL_LH_META_TRAFFIC_CLASS_NBITS-1
`define IRL_LH_META_TRAFFIC_CLASS `IRL_LH_META_TRAFFIC_CLASS_POS:0
`define IRL_LH_META_HDR_LEN_RANGE `IRL_LH_META_HDR_LEN_NBITS-1:0
`define IRL_LH_META_HDR_LEN_POS `IRL_LH_META_HDR_LEN_NBITS+`IRL_LH_META_TRAFFIC_CLASS_POS
`define IRL_LH_META_HDR_LEN `IRL_LH_META_HDR_LEN_POS:`IRL_LH_META_TRAFFIC_CLASS_POS+1
`define IRL_LH_META_BUF_PTR_RANGE `IRL_LH_META_BUF_PTR_NBITS-1:0
`define IRL_LH_META_BUF_PTR_POS `IRL_LH_META_BUF_PTR_NBITS+`IRL_LH_META_HDR_LEN_POS
`define IRL_LH_META_BUF_PTR `IRL_LH_META_BUF_PTR_POS:`IRL_LH_META_HDR_LEN_POS+1
`define IRL_LH_META_LEN_RANGE `IRL_LH_META_LEN_NBITS-1:0
`define IRL_LH_META_LEN_POS `IRL_LH_META_LEN_NBITS+`IRL_LH_META_BUF_PTR_POS
`define IRL_LH_META_LEN `IRL_LH_META_LEN_POS:`IRL_LH_META_BUF_PTR_POS+1
`define IRL_LH_META_PORT_RANGE `IRL_LH_META_PORT_NBITS-1:0
`define IRL_LH_META_PORT_POS `IRL_LH_META_PORT_NBITS+`IRL_LH_META_LEN_POS
`define IRL_LH_META_PORT `IRL_LH_META_PORT_POS:`IRL_LH_META_LEN_POS+1
`define IRL_LH_META_RCI_RANGE `IRL_LH_META_RCI_NBITS-1:0
`define IRL_LH_META_RCI_POS `IRL_LH_META_RCI_NBITS+`IRL_LH_META_PORT_POS
`define IRL_LH_META_RCI `IRL_LH_META_RCI_POS:`IRL_LH_META_PORT_POS+1
`define IRL_LH_META_FID_RANGE `IRL_LH_META_FID_NBITS-1:0
`define IRL_LH_META_FID_POS `IRL_LH_META_FID_NBITS+`IRL_LH_META_RCI_POS
`define IRL_LH_META_FID `IRL_LH_META_FID_POS:`IRL_LH_META_RCI_POS+1
`define IRL_LH_META_TID_RANGE `IRL_LH_META_TID_NBITS-1:0
`define IRL_LH_META_TID_POS `IRL_LH_META_TID_NBITS+`IRL_LH_META_FID_POS
`define IRL_LH_META_TID `IRL_LH_META_TID_POS:`IRL_LH_META_FID_POS+1
`define IRL_LH_META_TYPE1_RANGE `IRL_LH_META_TYPE1_NBITS-1:0
`define IRL_LH_META_TYPE1_POS `IRL_LH_META_TYPE1_NBITS+`IRL_LH_META_TID_POS
`define IRL_LH_META_TYPE1 `IRL_LH_META_TYPE1_POS:`IRL_LH_META_TID_POS+1
`define IRL_LH_META_TYPE3_RANGE `IRL_LH_META_TYPE3_NBITS-1:0
`define IRL_LH_META_TYPE3_POS `IRL_LH_META_TYPE3_NBITS+`IRL_LH_META_TYPE1_POS
`define IRL_LH_META_TYPE3 `IRL_LH_META_TYPE3_POS:`IRL_LH_META_TYPE1_POS+1
`define IRL_LH_META_DISCARD_RANGE `IRL_LH_META_DISCARD_NBITS-1:0
`define IRL_LH_META_DISCARD_POS `IRL_LH_META_DISCARD_NBITS+`IRL_LH_META_TYPE3_POS
`define IRL_LH_META_DISCARD `IRL_LH_META_DISCARD_POS:`IRL_LH_META_TYPE3_POS+1

`define LH_PP_META_HDR_LEN_NBITS `HEADER_LENGTH_NBITS
`define LH_PP_META_BUF_PTR_NBITS `BUF_PTR_NBITS
`define LH_PP_META_LEN_NBITS `PACKET_LENGTH_NBITS
`define LH_PP_META_PORT_NBITS `PORT_ID_NBITS
`define LH_PP_META_RCI_NBITS `RCI_NBITS
`define LH_PP_META_FID_NBITS `FID_NBITS
`define LH_PP_META_TID_NBITS `TID_NBITS
`define LH_PP_META_TYPE1_NBITS 1
`define LH_PP_META_TYPE3_NBITS 1
`define LH_PP_META_DISCARD_NBITS 1
`define LH_PP_META_NBITS `LH_PP_META_LEN_NBITS+`LH_PP_META_BUF_PTR_NBITS+`LH_PP_META_HDR_LEN_NBITS+`LH_PP_META_PORT_NBITS+`LH_PP_META_RCI_NBITS+`LH_PP_META_FID_NBITS+`LH_PP_META_TID_NBITS+`LH_PP_META_TYPE1_NBITS+`LH_PP_META_TYPE3_NBITS+`LH_PP_META_DISCARD_NBITS
`define LH_PP_META_RANGE `LH_PP_META_NBITS-1:0
`define LH_PP_META_HDR_LEN_RANGE `LH_PP_META_HDR_LEN_NBITS-1:0
`define LH_PP_META_HDR_LEN_POS `LH_PP_META_HDR_LEN_NBITS-1
`define LH_PP_META_HDR_LEN `LH_PP_META_HDR_LEN_POS:0
`define LH_PP_META_BUF_PTR_RANGE `LH_PP_META_BUF_PTR_NBITS-1:0
`define LH_PP_META_BUF_PTR_POS `LH_PP_META_BUF_PTR_NBITS+`LH_PP_META_HDR_LEN_POS
`define LH_PP_META_BUF_PTR `LH_PP_META_BUF_PTR_POS:`LH_PP_META_HDR_LEN_POS+1
`define LH_PP_META_LEN_RANGE `LH_PP_META_LEN_NBITS-1:0
`define LH_PP_META_LEN_POS `LH_PP_META_LEN_NBITS+`LH_PP_META_BUF_PTR_POS
`define LH_PP_META_LEN `LH_PP_META_LEN_POS:`LH_PP_META_BUF_PTR_POS+1
`define LH_PP_META_PORT_RANGE `LH_PP_META_PORT_NBITS-1:0
`define LH_PP_META_PORT_POS `LH_PP_META_PORT_NBITS+`LH_PP_META_LEN_POS
`define LH_PP_META_PORT `LH_PP_META_PORT_POS:`LH_PP_META_LEN_POS+1
`define LH_PP_META_RCI_RANGE `LH_PP_META_RCI_NBITS-1:0
`define LH_PP_META_RCI_POS `LH_PP_META_RCI_NBITS+`LH_PP_META_PORT_POS
`define LH_PP_META_RCI `LH_PP_META_RCI_POS:`LH_PP_META_PORT_POS+1
`define LH_PP_META_FID_RANGE `LH_PP_META_FID_NBITS-1:0
`define LH_PP_META_FID_POS `LH_PP_META_FID_NBITS+`LH_PP_META_RCI_POS
`define LH_PP_META_FID `LH_PP_META_FID_POS:`LH_PP_META_RCI_POS+1
`define LH_PP_META_TID_RANGE `LH_PP_META_TID_NBITS-1:0
`define LH_PP_META_TID_POS `LH_PP_META_TID_NBITS+`LH_PP_META_FID_POS
`define LH_PP_META_TID `LH_PP_META_TID_POS:`LH_PP_META_FID_POS+1
`define LH_PP_META_TYPE1_RANGE `LH_PP_META_TYPE1_NBITS-1:0
`define LH_PP_META_TYPE1_POS `LH_PP_META_TYPE1_NBITS+`LH_PP_META_TID_POS
`define LH_PP_META_TYPE1 `LH_PP_META_TYPE1_POS:`LH_PP_META_TID_POS+1
`define LH_PP_META_TYPE3_RANGE `LH_PP_META_TYPE3_NBITS-1:0
`define LH_PP_META_TYPE3_POS `LH_PP_META_TYPE3_NBITS+`LH_PP_META_TYPE1_POS
`define LH_PP_META_TYPE3 `LH_PP_META_TYPE3_POS:`LH_PP_META_TYPE1_POS+1
`define LH_PP_META_DISCARD_RANGE `LH_PP_META_DISCARD_NBITS-1:0
`define LH_PP_META_DISCARD_POS `LH_PP_META_DISCARD_NBITS+`LH_PP_META_TYPE3_POS
`define LH_PP_META_DISCARD `LH_PP_META_DISCARD_POS:`LH_PP_META_TYPE3_POS+1

`define LH_ECDSA_META_TRAFFIC_CLASS_NBITS `TRAFFIC_CLASS_NBITS
`define LH_ECDSA_META_HDR_LEN_NBITS `HEADER_LENGTH_NBITS
`define LH_ECDSA_META_BUF_PTR_NBITS `BUF_PTR_NBITS
`define LH_ECDSA_META_LEN_NBITS `PACKET_LENGTH_NBITS
`define LH_ECDSA_META_PORT_NBITS `PORT_ID_NBITS
`define LH_ECDSA_META_RCI_NBITS `RCI_NBITS
`define LH_ECDSA_META_FID_NBITS `FID_NBITS
`define LH_ECDSA_META_TID_NBITS `TID_NBITS
`define LH_ECDSA_META_TYPE1_NBITS 1
`define LH_ECDSA_META_TYPE3_NBITS 1
`define LH_ECDSA_META_DISCARD_NBITS 1
`define LH_ECDSA_META_NBITS `LH_ECDSA_META_TRAFFIC_CLASS_NBITS+`LH_ECDSA_META_LEN_NBITS+`LH_ECDSA_META_BUF_PTR_NBITS+`LH_ECDSA_META_HDR_LEN_NBITS+`LH_ECDSA_META_PORT_NBITS+`LH_ECDSA_META_RCI_NBITS+`LH_ECDSA_META_FID_NBITS+`LH_ECDSA_META_TID_NBITS+`LH_ECDSA_META_TYPE1_NBITS+`LH_ECDSA_META_TYPE3_NBITS+`LH_ECDSA_META_DISCARD_NBITS
`define LH_ECDSA_META_RANGE `LH_ECDSA_META_NBITS-1:0
`define LH_ECDSA_META_TRAFFIC_CLASS_RANGE `LH_ECDSA_META_TRAFFIC_CLASS_NBITS-1:0
`define LH_ECDSA_META_TRAFFIC_CLASS_POS `LH_ECDSA_META_TRAFFIC_CLASS_NBITS-1
`define LH_ECDSA_META_TRAFFIC_CLASS `LH_ECDSA_META_TRAFFIC_CLASS_POS:0
`define LH_ECDSA_META_HDR_LEN_RANGE `LH_ECDSA_META_HDR_LEN_NBITS-1:0
`define LH_ECDSA_META_HDR_LEN_POS `LH_ECDSA_META_HDR_LEN_NBITS+`LH_ECDSA_META_TRAFFIC_CLASS_POS
`define LH_ECDSA_META_HDR_LEN `LH_ECDSA_META_HDR_LEN_POS:`LH_ECDSA_META_TRAFFIC_CLASS_POS+1
`define LH_ECDSA_META_BUF_PTR_RANGE `LH_ECDSA_META_BUF_PTR_NBITS-1:0
`define LH_ECDSA_META_BUF_PTR_POS `LH_ECDSA_META_BUF_PTR_NBITS+`LH_ECDSA_META_HDR_LEN_POS
`define LH_ECDSA_META_BUF_PTR `LH_ECDSA_META_BUF_PTR_POS:`LH_ECDSA_META_HDR_LEN_POS+1
`define LH_ECDSA_META_LEN_RANGE `LH_ECDSA_META_LEN_NBITS-1:0
`define LH_ECDSA_META_LEN_POS `LH_ECDSA_META_LEN_NBITS+`LH_ECDSA_META_BUF_PTR_POS
`define LH_ECDSA_META_LEN `LH_ECDSA_META_LEN_POS:`LH_ECDSA_META_BUF_PTR_POS+1
`define LH_ECDSA_META_PORT_RANGE `LH_ECDSA_META_PORT_NBITS-1:0
`define LH_ECDSA_META_PORT_POS `LH_ECDSA_META_PORT_NBITS+`LH_ECDSA_META_LEN_POS
`define LH_ECDSA_META_PORT `LH_ECDSA_META_PORT_POS:`LH_ECDSA_META_LEN_POS+1
`define LH_ECDSA_META_RCI_RANGE `LH_ECDSA_META_RCI_NBITS-1:0
`define LH_ECDSA_META_RCI_POS `LH_ECDSA_META_RCI_NBITS+`LH_ECDSA_META_PORT_POS
`define LH_ECDSA_META_RCI `LH_ECDSA_META_RCI_POS:`LH_ECDSA_META_PORT_POS+1
`define LH_ECDSA_META_FID_RANGE `LH_ECDSA_META_FID_NBITS-1:0
`define LH_ECDSA_META_FID_POS `LH_ECDSA_META_FID_NBITS+`LH_ECDSA_META_RCI_POS
`define LH_ECDSA_META_FID `LH_ECDSA_META_FID_POS:`LH_ECDSA_META_RCI_POS+1
`define LH_ECDSA_META_TID_RANGE `LH_ECDSA_META_TID_NBITS-1:0
`define LH_ECDSA_META_TID_POS `LH_ECDSA_META_TID_NBITS+`LH_ECDSA_META_FID_POS
`define LH_ECDSA_META_TID `LH_ECDSA_META_TID_POS:`LH_ECDSA_META_FID_POS+1
`define LH_ECDSA_META_TYPE1_RANGE `LH_ECDSA_META_TYPE1_NBITS-1:0
`define LH_ECDSA_META_TYPE1_POS `LH_ECDSA_META_TYPE1_NBITS+`LH_ECDSA_META_TID_POS
`define LH_ECDSA_META_TYPE1 `LH_ECDSA_META_TYPE1_POS:`LH_ECDSA_META_TID_POS+1
`define LH_ECDSA_META_TYPE3_RANGE `LH_ECDSA_META_TYPE3_NBITS-1:0
`define LH_ECDSA_META_TYPE3_POS `LH_ECDSA_META_TYPE3_NBITS+`LH_ECDSA_META_TYPE1_POS
`define LH_ECDSA_META_TYPE3 `LH_ECDSA_META_TYPE3_POS:`LH_ECDSA_META_TYPE1_POS+1
`define LH_ECDSA_META_DISCARD_RANGE `LH_ECDSA_META_DISCARD_NBITS-1:0
`define LH_ECDSA_META_DISCARD_POS `LH_ECDSA_META_DISCARD_NBITS+`LH_ECDSA_META_TYPE3_POS
`define LH_ECDSA_META_DISCARD `LH_ECDSA_META_DISCARD_POS:`LH_ECDSA_META_TYPE3_POS+1

`define ECDSA_PP_META_DOMAIN_ID_NBITS `DOMAIN_ID_NBITS
`define ECDSA_PP_META_HDR_LEN_NBITS `HEADER_LENGTH_NBITS
`define ECDSA_PP_META_BUF_PTR_NBITS `BUF_PTR_NBITS
`define ECDSA_PP_META_LEN_NBITS `PACKET_LENGTH_NBITS
`define ECDSA_PP_META_PORT_NBITS `PORT_ID_NBITS
`define ECDSA_PP_META_RCI_NBITS `RCI_NBITS
`define ECDSA_PP_META_FID_NBITS `FID_NBITS
`define ECDSA_PP_META_TID_NBITS `TID_NBITS
`define ECDSA_PP_META_TYPE1_NBITS 1
`define ECDSA_PP_META_TYPE3_NBITS 1
`define ECDSA_PP_META_DISCARD_NBITS 1
`define ECDSA_PP_META_NBITS `ECDSA_PP_META_DOMAIN_ID_NBITS+`ECDSA_PP_META_LEN_NBITS+`ECDSA_PP_META_BUF_PTR_NBITS+`ECDSA_PP_META_HDR_LEN_NBITS+`ECDSA_PP_META_PORT_NBITS+`ECDSA_PP_META_RCI_NBITS+`ECDSA_PP_META_FID_NBITS+`ECDSA_PP_META_TID_NBITS+`ECDSA_PP_META_TYPE1_NBITS+`ECDSA_PP_META_TYPE3_NBITS+`ECDSA_PP_META_DISCARD_NBITS
`define ECDSA_PP_META_RANGE `ECDSA_PP_META_NBITS-1:0
`define ECDSA_PP_META_DOMAIN_ID_RANGE `ECDSA_PP_META_DOMAIN_ID_NBITS-1:0
`define ECDSA_PP_META_DOMAIN_ID_POS `ECDSA_PP_META_DOMAIN_ID_NBITS-1
`define ECDSA_PP_META_DOMAIN_ID `ECDSA_PP_META_DOMAIN_ID_POS:0
`define ECDSA_PP_META_HDR_LEN_RANGE `ECDSA_PP_META_HDR_LEN_NBITS-1:0
`define ECDSA_PP_META_HDR_LEN_POS `ECDSA_PP_META_HDR_LEN_NBITS+`ECDSA_PP_META_DOMAIN_ID_POS
`define ECDSA_PP_META_HDR_LEN `ECDSA_PP_META_HDR_LEN_POS:`ECDSA_PP_META_DOMAIN_ID_POS+1
`define ECDSA_PP_META_BUF_PTR_RANGE `ECDSA_PP_META_BUF_PTR_NBITS-1:0
`define ECDSA_PP_META_BUF_PTR_POS `ECDSA_PP_META_BUF_PTR_NBITS+`ECDSA_PP_META_HDR_LEN_POS
`define ECDSA_PP_META_BUF_PTR `ECDSA_PP_META_BUF_PTR_POS:`ECDSA_PP_META_HDR_LEN_POS+1
`define ECDSA_PP_META_LEN_RANGE `ECDSA_PP_META_LEN_NBITS-1:0
`define ECDSA_PP_META_LEN_POS `ECDSA_PP_META_LEN_NBITS+`ECDSA_PP_META_BUF_PTR_POS
`define ECDSA_PP_META_LEN `ECDSA_PP_META_LEN_POS:`ECDSA_PP_META_BUF_PTR_POS+1
`define ECDSA_PP_META_PORT_RANGE `ECDSA_PP_META_PORT_NBITS-1:0
`define ECDSA_PP_META_PORT_POS `ECDSA_PP_META_PORT_NBITS+`ECDSA_PP_META_LEN_POS
`define ECDSA_PP_META_PORT `ECDSA_PP_META_PORT_POS:`ECDSA_PP_META_LEN_POS+1
`define ECDSA_PP_META_RCI_RANGE `ECDSA_PP_META_RCI_NBITS-1:0
`define ECDSA_PP_META_RCI_POS `ECDSA_PP_META_RCI_NBITS+`ECDSA_PP_META_PORT_POS
`define ECDSA_PP_META_RCI `ECDSA_PP_META_RCI_POS:`ECDSA_PP_META_PORT_POS+1
`define ECDSA_PP_META_FID_RANGE `ECDSA_PP_META_FID_NBITS-1:0
`define ECDSA_PP_META_FID_POS `ECDSA_PP_META_FID_NBITS+`ECDSA_PP_META_RCI_POS
`define ECDSA_PP_META_FID `ECDSA_PP_META_FID_POS:`ECDSA_PP_META_RCI_POS+1
`define ECDSA_PP_META_TID_RANGE `ECDSA_PP_META_TID_NBITS-1:0
`define ECDSA_PP_META_TID_POS `ECDSA_PP_META_TID_NBITS+`ECDSA_PP_META_FID_POS
`define ECDSA_PP_META_TID `ECDSA_PP_META_TID_POS:`ECDSA_PP_META_FID_POS+1
`define ECDSA_PP_META_TYPE1_RANGE `ECDSA_PP_META_TYPE1_NBITS-1:0
`define ECDSA_PP_META_TYPE1_POS `ECDSA_PP_META_TYPE1_NBITS+`ECDSA_PP_META_TID_POS
`define ECDSA_PP_META_TYPE1 `ECDSA_PP_META_TYPE1_POS:`ECDSA_PP_META_TID_POS+1
`define ECDSA_PP_META_TYPE3_RANGE `ECDSA_PP_META_TYPE3_NBITS-1:0
`define ECDSA_PP_META_TYPE3_POS `ECDSA_PP_META_TYPE3_NBITS+`ECDSA_PP_META_TYPE1_POS
`define ECDSA_PP_META_TYPE3 `ECDSA_PP_META_TYPE3_POS:`ECDSA_PP_META_TYPE1_POS+1
`define ECDSA_PP_META_DISCARD_RANGE `ECDSA_PP_META_DISCARD_NBITS-1:0
`define ECDSA_PP_META_DISCARD_POS `ECDSA_PP_META_DISCARD_NBITS+`ECDSA_PP_META_TYPE3_POS
`define ECDSA_PP_META_DISCARD `ECDSA_PP_META_DISCARD_POS:`ECDSA_PP_META_TYPE3_POS+1

`define HOP_INFO_RCI_NBITS `RCI_NBITS
`define HOP_INFO_TYPE_NBITS 3
`define HOP_INFO_PC_NBITS 8
`define HOP_INFO_FLAGS_NBITS 8
`define HOP_INFO_BYTE_POINTER_NBITS 16
`define HOP_INFO_NBITS `HOP_INFO_RCI_NBITS+`HOP_INFO_TYPE_NBITS+`HOP_INFO_PC_NBITS+`HOP_INFO_FLAGS_NBITS+`HOP_INFO_BYTE_POINTER_NBITS
`define HOP_INFO_RANGE `HOP_INFO_NBITS-1:0
`define HOP_INFO_RCI_RANGE `HOP_INFO_RCI_NBITS-1:0
`define HOP_INFO_RCI_POS `HOP_INFO_RCI_NBITS-1
`define HOP_INFO_RCI `HOP_INFO_RCI_POS:0
`define HOP_INFO_TYPE_RANGE `HOP_INFO_TYPE_NBITS-1:0
`define HOP_INFO_TYPE_POS `HOP_INFO_TYPE_NBITS+`HOP_INFO_RCI_POS
`define HOP_INFO_TYPE `HOP_INFO_TYPE_POS:`HOP_INFO_RCI_POS+1
`define HOP_INFO_PC_RANGE `HOP_INFO_PC_NBITS-1:0
`define HOP_INFO_PC_POS `HOP_INFO_PC_NBITS+`HOP_INFO_TYPE_POS
`define HOP_INFO_PC `HOP_INFO_PC_POS:`HOP_INFO_TYPE_POS+1
`define HOP_INFO_FLAGS_RANGE `HOP_INFO_FLAGS_NBITS-1:0
`define HOP_INFO_FLAGS_POS `HOP_INFO_FLAGS_NBITS+`HOP_INFO_PC_POS
`define HOP_INFO_FLAGS `HOP_INFO_FLAGS_POS:`HOP_INFO_PC_POS+1
`define HOP_INFO_BYTE_POINTER_RANGE `HOP_INFO_BYTE_POINTER_NBITS-1:0
`define HOP_INFO_BYTE_POINTER_POS `HOP_INFO_BYTE_POINTER_NBITS+`HOP_INFO_FLAGS_POS
`define HOP_INFO_BYTE_POINTER `HOP_INFO_BYTE_POINTER_POS:`HOP_INFO_FLAGS_POS+1

`define PU_HOP_META_TIME_NBITS 32
`define PU_HOP_META_RCI_NBITS 16
`define PU_HOP_META_PKT_TYPE_NBITS 8
`define PU_HOP_META_SWITCH_TAG_NBITS `SWITCH_TAG_NBITS
`define PU_HOP_META_F_PAYLOAD_NBITS `FLOW_PU_NBITS
`define PU_HOP_META_TID_NBITS `TID_NBITS
`define PU_HOP_META_FID_NBITS `FID_NBITS
`define PU_HOP_META_NBITS `PU_HOP_META_TIME_NBITS+`PU_HOP_META_SWITCH_TAG_NBITS+`PU_HOP_META_PKT_TYPE_NBITS+`PU_HOP_META_RCI_NBITS+`PU_HOP_META_F_PAYLOAD_NBITS+`PU_HOP_META_TID_NBITS+`PU_HOP_META_FID_NBITS
`define PU_HOP_META_RANGE `PU_HOP_META_NBITS-1:0
`define PU_HOP_META_TIME_RANGE `PU_HOP_META_TIME_NBITS-1:0
`define PU_HOP_META_TIME_POS `PU_HOP_META_TIME_NBITS-1
`define PU_HOP_META_TIME `PU_HOP_META_TIME_POS:0
`define PU_HOP_META_RCI_RANGE `PU_HOP_META_RCI_NBITS-1:0
`define PU_HOP_META_RCI_POS `PU_HOP_META_RCI_NBITS+`PU_HOP_META_TIME_POS
`define PU_HOP_META_RCI `PU_HOP_META_RCI_POS:`PU_HOP_META_TIME_POS+1
`define PU_HOP_META_PKT_TYPE_RANGE `PU_HOP_META_PKT_TYPE_NBITS-1:0
`define PU_HOP_META_PKT_TYPE_POS `PU_HOP_META_PKT_TYPE_NBITS+`PU_HOP_META_RCI_POS
`define PU_HOP_META_PKT_TYPE `PU_HOP_META_PKT_TYPE_POS:`PU_HOP_META_RCI_POS+1
`define PU_HOP_META_SWITCH_TAG_RANGE `PU_HOP_META_SWITCH_TAG_NBITS-1:0
`define PU_HOP_META_SWITCH_TAG_POS `PU_HOP_META_SWITCH_TAG_NBITS+`PU_HOP_META_PKT_TYPE_POS
`define PU_HOP_META_SWITCH_TAG `PU_HOP_META_SWITCH_TAG_POS:`PU_HOP_META_PKT_TYPE_POS+1
`define PU_HOP_META_F_PAYLOAD_RANGE `PU_HOP_META_F_PAYLOAD_NBITS-1:0
`define PU_HOP_META_F_PAYLOAD_POS `PU_HOP_META_F_PAYLOAD_NBITS+`PU_HOP_META_SWITCH_TAG_POS
`define PU_HOP_META_F_PAYLOAD `PU_HOP_META_F_PAYLOAD_POS:`PU_HOP_META_SWITCH_TAG_POS+1
`define PU_HOP_META_TID_RANGE `PU_HOP_META_TID_NBITS-1:0
`define PU_HOP_META_TID_POS `PU_HOP_META_TID_NBITS+`PU_HOP_META_F_PAYLOAD_POS
`define PU_HOP_META_TID `PU_HOP_META_TID_POS:`PU_HOP_META_F_PAYLOAD_POS+1
`define PU_HOP_META_FID_RANGE `PU_HOP_META_FID_NBITS-1:0
`define PU_HOP_META_FID_POS `PU_HOP_META_FID_NBITS+`PU_HOP_META_TID_POS
`define PU_HOP_META_FID `PU_HOP_META_FID_POS:`PU_HOP_META_TID_POS+1

`define ENQ_ED_CMD_PTR_UPDATE_NBITS 1
`define ENQ_ED_CMD_CUR_PTR_NBITS 16
`define ENQ_ED_CMD_PTR_LOC_NBITS 10
`define ENQ_ED_CMD_PD_UPDATE_NBITS 1
`define ENQ_ED_CMD_PD_LEN_NBITS 7
`define ENQ_ED_CMD_PD_LOC_NBITS 10
`define ENQ_ED_CMD_PD_BP_NBITS 10
`define ENQ_ED_CMD_OUT_RCI_NBITS `RCI_NBITS
`define ENQ_ED_CMD_PKT_LEN_NBITS `PACKET_LENGTH_NBITS
`define ENQ_ED_CMD_NBITS `ENQ_ED_CMD_PKT_LEN_NBITS+`ENQ_ED_CMD_OUT_RCI_NBITS+`ENQ_ED_CMD_PD_BP_NBITS+`ENQ_ED_CMD_PD_LOC_NBITS+`ENQ_ED_CMD_PD_LEN_NBITS+`ENQ_ED_CMD_PD_UPDATE_NBITS+`ENQ_ED_CMD_PTR_LOC_NBITS+`ENQ_ED_CMD_CUR_PTR_NBITS+`ENQ_ED_CMD_PTR_UPDATE_NBITS
`define ENQ_ED_CMD_RANGE `ENQ_ED_CMD_NBITS-1:0
`define ENQ_ED_CMD_PTR_UPDATE_RANGE `ENQ_ED_CMD_PTR_UPDATE_NBITS-1:0
`define ENQ_ED_CMD_PTR_UPDATE_POS `ENQ_ED_CMD_PTR_UPDATE_NBITS-1
`define ENQ_ED_CMD_PTR_UPDATE `ENQ_ED_CMD_PTR_UPDATE_POS:0
`define ENQ_ED_CMD_CUR_PTR_RANGE `ENQ_ED_CMD_CUR_PTR_NBITS-1:0
`define ENQ_ED_CMD_CUR_PTR_POS `ENQ_ED_CMD_CUR_PTR_NBITS+`ENQ_ED_CMD_PTR_UPDATE_POS
`define ENQ_ED_CMD_CUR_PTR `ENQ_ED_CMD_CUR_PTR_POS:`ENQ_ED_CMD_PTR_UPDATE_POS+1
`define ENQ_ED_CMD_PTR_LOC_RANGE `ENQ_ED_CMD_PTR_LOC_NBITS-1:0
`define ENQ_ED_CMD_PTR_LOC_POS `ENQ_ED_CMD_PTR_LOC_NBITS+`ENQ_ED_CMD_CUR_PTR_POS
`define ENQ_ED_CMD_PTR_LOC `ENQ_ED_CMD_PTR_LOC_POS:`ENQ_ED_CMD_CUR_PTR_POS+1
`define ENQ_ED_CMD_PD_UPDATE_RANGE `ENQ_ED_CMD_PD_UPDATE_NBITS-1:0
`define ENQ_ED_CMD_PD_UPDATE_POS `ENQ_ED_CMD_PD_UPDATE_NBITS+`ENQ_ED_CMD_PTR_LOC_POS
`define ENQ_ED_CMD_PD_UPDATE `ENQ_ED_CMD_PD_UPDATE_POS:`ENQ_ED_CMD_PTR_LOC_POS+1
`define ENQ_ED_CMD_PD_LEN_RANGE `ENQ_ED_CMD_PD_LEN_NBITS-1:0
`define ENQ_ED_CMD_PD_LEN_POS `ENQ_ED_CMD_PD_LEN_NBITS+`ENQ_ED_CMD_PD_UPDATE_POS
`define ENQ_ED_CMD_PD_LEN `ENQ_ED_CMD_PD_LEN_POS:`ENQ_ED_CMD_PD_UPDATE_POS+1
`define ENQ_ED_CMD_PD_LOC_RANGE `ENQ_ED_CMD_PD_LOC_NBITS-1:0
`define ENQ_ED_CMD_PD_LOC_POS `ENQ_ED_CMD_PD_LOC_NBITS+`ENQ_ED_CMD_PD_LEN_POS
`define ENQ_ED_CMD_PD_LOC `ENQ_ED_CMD_PD_LOC_POS:`ENQ_ED_CMD_PD_LEN_POS+1
`define ENQ_ED_CMD_PD_BP_RANGE `ENQ_ED_CMD_PD_BP_NBITS-1:0
`define ENQ_ED_CMD_PD_BP_POS `ENQ_ED_CMD_PD_BP_NBITS+`ENQ_ED_CMD_PD_LOC_POS
`define ENQ_ED_CMD_PD_BP `ENQ_ED_CMD_PD_BP_POS:`ENQ_ED_CMD_PD_LOC_POS+1
`define ENQ_ED_CMD_OUT_RCI_RANGE `ENQ_ED_CMD_OUT_RCI_NBITS-1:0
`define ENQ_ED_CMD_OUT_RCI_POS `ENQ_ED_CMD_OUT_RCI_NBITS+`ENQ_ED_CMD_PD_BP_POS
`define ENQ_ED_CMD_OUT_RCI `ENQ_ED_CMD_OUT_RCI_POS:`ENQ_ED_CMD_PD_BP_POS+1
`define ENQ_ED_CMD_PKT_LEN_RANGE `ENQ_ED_CMD_PKT_LEN_NBITS-1:0
`define ENQ_ED_CMD_PKT_LEN_POS `ENQ_ED_CMD_PKT_LEN_NBITS+`ENQ_ED_CMD_OUT_RCI_POS
`define ENQ_ED_CMD_PKT_LEN `ENQ_ED_CMD_PKT_LEN_POS:`ENQ_ED_CMD_OUT_RCI_POS+1

`define ENQ_ED_CMD_PTR_LOC_NBITS 10
`define ENQ_ED_CMD_PD_LOC_NBITS 10

`define PP_PIARB_META_PTR_LOC_NBITS `ENQ_ED_CMD_PTR_LOC_NBITS
`define PP_PIARB_META_PD_LOC_NBITS `ENQ_ED_CMD_PD_LOC_NBITS
`define PP_PIARB_META_DOMAIN_ID_NBITS `DOMAIN_ID_NBITS
`define PP_PIARB_META_HDR_LEN_NBITS `HEADER_LENGTH_NBITS
`define PP_PIARB_META_BUF_PTR_NBITS `BUF_PTR_NBITS
`define PP_PIARB_META_LEN_NBITS `PACKET_LENGTH_NBITS
`define PP_PIARB_META_PORT_NBITS `PORT_ID_NBITS
`define PP_PIARB_META_RCI_NBITS `RCI_NBITS
`define PP_PIARB_META_FID_SEL_NBITS 1
`define PP_PIARB_META_FID_NBITS `FID_NBITS
`define PP_PIARB_META_TID_NBITS `TID_NBITS
`define PP_PIARB_META_TYPE1_NBITS 1
`define PP_PIARB_META_TYPE3_NBITS 1
`define PP_PIARB_META_TIME_NBITS 32
`define PP_PIARB_META_DISCARD_NBITS 1
`define PP_PIARB_META_NBITS `PP_PIARB_META_PTR_LOC_NBITS+`PP_PIARB_META_PD_LOC_NBITS+`PP_PIARB_META_DOMAIN_ID_NBITS+`PP_PIARB_META_LEN_NBITS+`PP_PIARB_META_BUF_PTR_NBITS+`PP_PIARB_META_HDR_LEN_NBITS+`PP_PIARB_META_PORT_NBITS+`PP_PIARB_META_RCI_NBITS+`PP_PIARB_META_FID_SEL_NBITS+`PP_PIARB_META_FID_NBITS+`PP_PIARB_META_TID_NBITS+`PP_PIARB_META_TYPE1_NBITS+`PP_PIARB_META_TYPE3_NBITS+`PP_PIARB_META_TIME_NBITS+`PP_PIARB_META_DISCARD_NBITS
`define PP_PIARB_META_RANGE `PP_PIARB_META_NBITS-1:0
`define PP_PIARB_META_PTR_LOC_RANGE `PP_PIARB_META_PTR_LOC_NBITS-1:0
`define PP_PIARB_META_PTR_LOC_POS `PP_PIARB_META_PTR_LOC_NBITS-1
`define PP_PIARB_META_PTR_LOC `PP_PIARB_META_PTR_LOC_POS:0
`define PP_PIARB_META_PD_LOC_RANGE `PP_PIARB_META_PD_LOC_NBITS-1:0
`define PP_PIARB_META_PD_LOC_POS `PP_PIARB_META_PD_LOC_NBITS+`PP_PIARB_META_PTR_LOC_POS
`define PP_PIARB_META_PD_LOC `PP_PIARB_META_PD_LOC_POS:PP_PIARB_META_PTR_LOC_POS+1
`define PP_PIARB_META_DOMAIN_ID_RANGE `PP_PIARB_META_DOMAIN_ID_NBITS-1:0
`define PP_PIARB_META_DOMAIN_ID_POS `PP_PIARB_META_DOMAIN_ID_NBITS+`PP_PIARB_META_PD_LOC_POS
`define PP_PIARB_META_DOMAIN_ID `PP_PIARB_META_DOMAIN_ID_POS:PP_PIARB_META_PD_LOC_POS+1
`define PP_PIARB_META_HDR_LEN_RANGE `PP_PIARB_META_HDR_LEN_NBITS-1:0
`define PP_PIARB_META_HDR_LEN_POS `PP_PIARB_META_HDR_LEN_NBITS+`PP_PIARB_META_DOMAIN_ID_POS
`define PP_PIARB_META_HDR_LEN `PP_PIARB_META_HDR_LEN_POS:PP_PIARB_META_DOMAIN_ID_POS+1
`define PP_PIARB_META_BUF_PTR_RANGE `PP_PIARB_META_BUF_PTR_NBITS-1:0
`define PP_PIARB_META_BUF_PTR_POS `PP_PIARB_META_BUF_PTR_NBITS+`PP_PIARB_META_HDR_LEN_POS
`define PP_PIARB_META_BUF_PTR `PP_PIARB_META_BUF_PTR_POS:`PP_PIARB_META_HDR_LEN_POS+1
`define PP_PIARB_META_LEN_RANGE `PP_PIARB_META_LEN_NBITS-1:0
`define PP_PIARB_META_LEN_POS `PP_PIARB_META_LEN_NBITS+`PP_PIARB_META_BUF_PTR_POS
`define PP_PIARB_META_LEN `PP_PIARB_META_LEN_POS:`PP_PIARB_META_BUF_PTR_POS+1
`define PP_PIARB_META_PORT_RANGE `PP_PIARB_META_PORT_NBITS-1:0
`define PP_PIARB_META_PORT_POS `PP_PIARB_META_PORT_NBITS+`PP_PIARB_META_LEN_POS
`define PP_PIARB_META_PORT `PP_PIARB_META_PORT_POS:`PP_PIARB_META_LEN_POS+1
`define PP_PIARB_META_RCI_RANGE `PP_PIARB_META_RCI_NBITS-1:0
`define PP_PIARB_META_RCI_POS `PP_PIARB_META_RCI_NBITS+`PP_PIARB_META_PORT_POS
`define PP_PIARB_META_RCI `PP_PIARB_META_RCI_POS:`PP_PIARB_META_PORT_POS+1
`define PP_PIARB_META_FID_SEL_RANGE `PP_PIARB_META_FID_SEL_NBITS-1:0
`define PP_PIARB_META_FID_SEL_POS `PP_PIARB_META_FID_SEL_NBITS+`PP_PIARB_META_RCI_POS
`define PP_PIARB_META_FID_SEL `PP_PIARB_META_FID_SEL_POS:`PP_PIARB_META_RCI_POS+1
`define PP_PIARB_META_FID_RANGE `PP_PIARB_META_FID_NBITS-1:0
`define PP_PIARB_META_FID_POS `PP_PIARB_META_FID_NBITS+`PP_PIARB_META_FID_SEL_POS
`define PP_PIARB_META_FID `PP_PIARB_META_FID_POS:`PP_PIARB_META_FID_SEL_POS+1
`define PP_PIARB_META_TID_RANGE `PP_PIARB_META_TID_NBITS-1:0
`define PP_PIARB_META_TID_POS `PP_PIARB_META_TID_NBITS+`PP_PIARB_META_FID_POS
`define PP_PIARB_META_TID `PP_PIARB_META_TID_POS:`PP_PIARB_META_FID_POS+1
`define PP_PIARB_META_TYPE1_RANGE `PP_PIARB_META_TYPE1_NBITS-1:0
`define PP_PIARB_META_TYPE1_POS `PP_PIARB_META_TYPE1_NBITS+`PP_PIARB_META_TID_POS
`define PP_PIARB_META_TYPE1 `PP_PIARB_META_TYPE1_POS:`PP_PIARB_META_TID_POS+1
`define PP_PIARB_META_TYPE3_RANGE `PP_PIARB_META_TYPE3_NBITS-1:0
`define PP_PIARB_META_TYPE3_POS `PP_PIARB_META_TYPE3_NBITS+`PP_PIARB_META_TYPE1_POS
`define PP_PIARB_META_TYPE3 `PP_PIARB_META_TYPE3_POS:`PP_PIARB_META_TYPE1_POS+1
`define PP_PIARB_META_TIME_RANGE `PP_PIARB_META_TIME_NBITS-1:0
`define PP_PIARB_META_TIME_POS `PP_PIARB_META_TIME_NBITS+`PP_PIARB_META_TYPE3_POS
`define PP_PIARB_META_TIME `PP_PIARB_META_TIME_POS:`PP_PIARB_META_TYPE3_POS+1
`define PP_PIARB_META_DISCARD_RANGE `PP_PIARB_META_DISCARD_NBITS-1:0
`define PP_PIARB_META_DISCARD_POS `PP_PIARB_META_DISCARD_NBITS+`PP_PIARB_META_TIME_POS
`define PP_PIARB_META_DISCARD `PP_PIARB_META_DISCARD_POS:`PP_PIARB_META_TIME_POS+1

`define PIARB_ASA_META_DOMAIN_ID_NBITS `DOMAIN_ID_NBITS
`define PIARB_ASA_META_HDR_LEN_NBITS `HEADER_LENGTH_NBITS
`define PIARB_ASA_META_BUF_PTR_NBITS `BUF_PTR_NBITS
`define PIARB_ASA_META_LEN_NBITS `PACKET_LENGTH_NBITS
`define PIARB_ASA_META_PORT_NBITS `PORT_ID_NBITS
`define PIARB_ASA_META_RCI_NBITS `RCI_NBITS
`define PIARB_ASA_META_FID_SEL_NBITS 1
`define PIARB_ASA_META_FID_NBITS `FID_NBITS
`define PIARB_ASA_META_TID_NBITS `TID_NBITS
`define PIARB_ASA_META_TYPE1_NBITS 1
`define PIARB_ASA_META_TYPE3_NBITS 1
`define PIARB_ASA_META_TIME_NBITS 32
`define PIARB_ASA_META_DISCARD_NBITS 1
`define PIARB_ASA_META_NBITS `PIARB_ASA_META_DOMAIN_ID_NBITS+`PIARB_ASA_META_LEN_NBITS+`PIARB_ASA_META_BUF_PTR_NBITS+`PIARB_ASA_META_HDR_LEN_NBITS+`PIARB_ASA_META_PORT_NBITS+`PIARB_ASA_META_RCI_NBITS+`PIARB_ASA_META_FID_SEL_NBITS+`PIARB_ASA_META_FID_NBITS+`PIARB_ASA_META_TID_NBITS+`PIARB_ASA_META_TYPE1_NBITS+`PIARB_ASA_META_TYPE3_NBITS+`PIARB_ASA_META_TIME_NBITS+`PIARB_ASA_META_DISCARD_NBITS
`define PIARB_ASA_META_RANGE `PIARB_ASA_META_NBITS-1:0
`define PIARB_ASA_META_DOMAIN_ID_RANGE `PIARB_ASA_META_DOMAIN_ID_NBITS-1:0
`define PIARB_ASA_META_DOMAIN_ID_POS `PIARB_ASA_META_DOMAIN_ID_NBITS-1
`define PIARB_ASA_META_DOMAIN_ID `PIARB_ASA_META_DOMAIN_ID_POS:0
`define PIARB_ASA_META_HDR_LEN_RANGE `PIARB_ASA_META_HDR_LEN_NBITS-1:0
`define PIARB_ASA_META_HDR_LEN_POS `PIARB_ASA_META_HDR_LEN_NBITS+`PIARB_ASA_META_DOMAIN_ID_POS
`define PIARB_ASA_META_HDR_LEN `PIARB_ASA_META_HDR_LEN_POS:PIARB_ASA_META_DOMAIN_ID_POS+1
`define PIARB_ASA_META_BUF_PTR_RANGE `PIARB_ASA_META_BUF_PTR_NBITS-1:0
`define PIARB_ASA_META_BUF_PTR_POS `PIARB_ASA_META_BUF_PTR_NBITS+`PIARB_ASA_META_HDR_LEN_POS
`define PIARB_ASA_META_BUF_PTR `PIARB_ASA_META_BUF_PTR_POS:`PIARB_ASA_META_HDR_LEN_POS+1
`define PIARB_ASA_META_LEN_RANGE `PIARB_ASA_META_LEN_NBITS-1:0
`define PIARB_ASA_META_LEN_POS `PIARB_ASA_META_LEN_NBITS+`PIARB_ASA_META_BUF_PTR_POS
`define PIARB_ASA_META_LEN `PIARB_ASA_META_LEN_POS:`PIARB_ASA_META_BUF_PTR_POS+1
`define PIARB_ASA_META_PORT_RANGE `PIARB_ASA_META_PORT_NBITS-1:0
`define PIARB_ASA_META_PORT_POS `PIARB_ASA_META_PORT_NBITS+`PIARB_ASA_META_LEN_POS
`define PIARB_ASA_META_PORT `PIARB_ASA_META_PORT_POS:`PIARB_ASA_META_LEN_POS+1
`define PIARB_ASA_META_RCI_RANGE `PIARB_ASA_META_RCI_NBITS-1:0
`define PIARB_ASA_META_RCI_POS `PIARB_ASA_META_RCI_NBITS+`PIARB_ASA_META_PORT_POS
`define PIARB_ASA_META_RCI `PIARB_ASA_META_RCI_POS:`PIARB_ASA_META_PORT_POS+1
`define PIARB_ASA_META_FID_SEL_RANGE `PIARB_ASA_META_FID_SEL_NBITS-1:0
`define PIARB_ASA_META_FID_SEL_POS `PIARB_ASA_META_FID_SEL_NBITS+`PIARB_ASA_META_RCI_POS
`define PIARB_ASA_META_FID_SEL `PIARB_ASA_META_FID_SEL_POS:`PIARB_ASA_META_RCI_POS+1
`define PIARB_ASA_META_FID_RANGE `PIARB_ASA_META_FID_NBITS-1:0
`define PIARB_ASA_META_FID_POS `PIARB_ASA_META_FID_NBITS+`PIARB_ASA_META_FID_SEL_POS
`define PIARB_ASA_META_FID `PIARB_ASA_META_FID_POS:`PIARB_ASA_META_FID_SEL_POS+1
`define PIARB_ASA_META_TID_RANGE `PIARB_ASA_META_TID_NBITS-1:0
`define PIARB_ASA_META_TID_POS `PIARB_ASA_META_TID_NBITS+`PIARB_ASA_META_FID_POS
`define PIARB_ASA_META_TID `PIARB_ASA_META_TID_POS:`PIARB_ASA_META_FID_POS+1
`define PIARB_ASA_META_TYPE1_RANGE `PIARB_ASA_META_TYPE1_NBITS-1:0
`define PIARB_ASA_META_TYPE1_POS `PIARB_ASA_META_TYPE1_NBITS+`PIARB_ASA_META_TID_POS
`define PIARB_ASA_META_TYPE1 `PIARB_ASA_META_TYPE1_POS:`PIARB_ASA_META_TID_POS+1
`define PIARB_ASA_META_TYPE3_RANGE `PIARB_ASA_META_TYPE3_NBITS-1:0
`define PIARB_ASA_META_TYPE3_POS `PIARB_ASA_META_TYPE3_NBITS+`PIARB_ASA_META_TYPE1_POS
`define PIARB_ASA_META_TYPE3 `PIARB_ASA_META_TYPE3_POS:`PIARB_ASA_META_TYPE1_POS+1
`define PIARB_ASA_META_TIME_RANGE `PIARB_ASA_META_TIME_NBITS-1:0
`define PIARB_ASA_META_TIME_POS `PIARB_ASA_META_TIME_NBITS+`PIARB_ASA_META_TYPE3_POS
`define PIARB_ASA_META_TIME `PIARB_ASA_META_TIME_POS:`PIARB_ASA_META_TYPE3_POS+1
`define PIARB_ASA_META_DISCARD_RANGE `PIARB_ASA_META_DISCARD_NBITS-1:0
`define PIARB_ASA_META_DISCARD_POS `PIARB_ASA_META_DISCARD_NBITS+`PIARB_ASA_META_TIME_POS
`define PIARB_ASA_META_DISCARD `PIARB_ASA_META_DISCARD_POS:`PIARB_ASA_META_TIME_POS+1

`define PP_META_DOMAIN_ID_NBITS `DOMAIN_ID_NBITS
`define PP_META_HDR_LEN_NBITS `HEADER_LENGTH_NBITS
`define PP_META_BUF_PTR_NBITS `BUF_PTR_NBITS
`define PP_META_LEN_NBITS `PACKET_LENGTH_NBITS
`define PP_META_PORT_NBITS `PORT_ID_NBITS
`define PP_META_RCI_NBITS `RCI_NBITS
`define PP_META_FID_SEL_NBITS 1
`define PP_META_FID_NBITS `FID_NBITS
`define PP_META_TID_NBITS `TID_NBITS
`define PP_META_TYPE1_NBITS 1
`define PP_META_TYPE3_NBITS 1
`define PP_META_DISCARD_NBITS 1
`define PP_META_NBITS `PP_META_DOMAIN_ID_NBITS+`PP_META_LEN_NBITS+`PP_META_BUF_PTR_NBITS+`PP_META_HDR_LEN_NBITS+`PP_META_PORT_NBITS+`PP_META_RCI_NBITS+`PP_META_FID_NBITS+`PP_META_TID_NBITS+`PP_META_TYPE1_NBITS+`PP_META_TYPE3_NBITS+`PP_META_DISCARD_NBITS
`define PP_META_RANGE `PP_META_NBITS-1:0
`define PP_META_DOMAIN_ID_RANGE `PP_META_DOMAIN_ID_NBITS-1:0
`define PP_META_DOMAIN_ID_POS `PP_META_DOMAIN_ID_NBITS-1
`define PP_META_DOMAIN_ID `PP_META_DOMAIN_ID_POS:0
`define PP_META_HDR_LEN_RANGE `PP_META_HDR_LEN_NBITS-1:0
`define PP_META_HDR_LEN_POS `PP_META_HDR_LEN_NBITS+`PP_META_DOMAIN_ID_POS
`define PP_META_HDR_LEN `PP_META_HDR_LEN_POS:PP_META_DOMAIN_ID_POS+1
`define PP_META_BUF_PTR_RANGE `PP_META_BUF_PTR_NBITS-1:0
`define PP_META_BUF_PTR_POS `PP_META_BUF_PTR_NBITS+`PP_META_HDR_LEN_POS
`define PP_META_BUF_PTR `PP_META_BUF_PTR_POS:`PP_META_HDR_LEN_POS+1
`define PP_META_LEN_RANGE `PP_META_LEN_NBITS-1:0
`define PP_META_LEN_POS `PP_META_LEN_NBITS+`PP_META_BUF_PTR_POS
`define PP_META_LEN `PP_META_LEN_POS:`PP_META_BUF_PTR_POS+1
`define PP_META_PORT_RANGE `PP_META_PORT_NBITS-1:0
`define PP_META_PORT_POS `PP_META_PORT_NBITS+`PP_META_LEN_POS
`define PP_META_PORT `PP_META_PORT_POS:`PP_META_LEN_POS+1
`define PP_META_RCI_RANGE `PP_META_RCI_NBITS-1:0
`define PP_META_RCI_POS `PP_META_RCI_NBITS+`PP_META_PORT_POS
`define PP_META_RCI `PP_META_RCI_POS:`PP_META_PORT_POS+1
`define PP_META_FID_RANGE `PP_META_FID_NBITS-1:0
`define PP_META_FID_POS `PP_META_FID_NBITS+`PP_META_RCI_POS
`define PP_META_FID `PP_META_FID_POS:`PP_META_RCI_POS+1
`define PP_META_TID_RANGE `PP_META_TID_NBITS-1:0
`define PP_META_TID_POS `PP_META_TID_NBITS+`PP_META_FID_POS
`define PP_META_TID `PP_META_TID_POS:`PP_META_FID_POS+1
`define PP_META_TYPE1_RANGE `PP_META_TYPE1_NBITS-1:0
`define PP_META_TYPE1_POS `PP_META_TYPE1_NBITS+`PP_META_TID_POS
`define PP_META_TYPE1 `PP_META_TYPE1_POS:`PP_META_TID_POS+1
`define PP_META_TYPE3_RANGE `PP_META_TYPE3_NBITS-1:0
`define PP_META_TYPE3_POS `PP_META_TYPE3_NBITS+`PP_META_TYPE1_POS
`define PP_META_TYPE3 `PP_META_TYPE3_POS:`PP_META_TYPE1_POS+1
`define PP_META_DISCARD_RANGE `PP_META_DISCARD_NBITS-1:0
`define PP_META_DISCARD_POS `PP_META_DISCARD_NBITS+`PP_META_TYPE3_POS
`define PP_META_DISCARD `PP_META_DISCARD_POS:`PP_META_TYPE3_POS+1

`define PP_PU_META_LEN_NBITS `PACKET_LENGTH_NBITS
`define PP_PU_META_PORT_NBITS `PORT_ID_NBITS
`define PP_PU_META_RCI_NBITS `RCI_NBITS
`define PP_PU_META_FID_NBITS `FID_NBITS
`define PP_PU_META_TID_NBITS `TID_NBITS
`define PP_PU_META_TYPE1_NBITS 1
`define PP_PU_META_F_PAYLOAD_NBITS `FLOW_PU_NBITS
`define PP_PU_META_T_PAYLOAD_NBITS `SWITCH_TAG_NBITS
`define PP_PU_META_NBITS `PP_PU_META_LEN_NBITS+`PP_PU_META_PORT_NBITS+`PP_PU_META_RCI_NBITS+`PP_PU_META_FID_NBITS+`PP_PU_META_TID_NBITS+`PP_PU_META_TYPE1_NBITS+`PP_PU_META_F_PAYLOAD_NBITS+`PP_PU_META_T_PAYLOAD_NBITS
`define PP_PU_META_RANGE `PP_PU_META_NBITS-1:0
`define PP_PU_META_LEN_RANGE `PP_PU_META_LEN_NBITS-1:0
`define PP_PU_META_LEN_POS `PP_PU_META_LEN_NBITS-1
`define PP_PU_META_LEN `PP_PU_META_LEN_POS:0
`define PP_PU_META_PORT_RANGE `PP_PU_META_PORT_NBITS-1:0
`define PP_PU_META_PORT_POS `PP_PU_META_PORT_NBITS+`PP_PU_META_LEN_POS
`define PP_PU_META_PORT `PP_PU_META_PORT_POS:`PP_PU_META_LEN_POS+1
`define PP_PU_META_RCI_RANGE `PP_PU_META_RCI_NBITS-1:0
`define PP_PU_META_RCI_POS `PP_PU_META_RCI_NBITS+`PP_PU_META_PORT_POS
`define PP_PU_META_RCI `PP_PU_META_RCI_POS:`PP_PU_META_PORT_POS+1
`define PP_PU_META_FID_RANGE `PP_PU_META_FID_NBITS-1:0
`define PP_PU_META_FID_POS `PP_PU_META_FID_NBITS+`PP_PU_META_RCI_POS
`define PP_PU_META_FID `PP_PU_META_FID_POS:`PP_PU_META_RCI_POS+1
`define PP_PU_META_TID_RANGE `PP_PU_META_TID_NBITS-1:0
`define PP_PU_META_TID_POS `PP_PU_META_TID_NBITS+`PP_PU_META_FID_POS
`define PP_PU_META_TID `PP_PU_META_TID_POS:`PP_PU_META_FID_POS+1
`define PP_PU_META_TYPE1_RANGE `PP_PU_META_TYPE1_NBITS-1:0
`define PP_PU_META_TYPE1_POS `PP_PU_META_TYPE1_NBITS+`PP_PU_META_TID_POS
`define PP_PU_META_TYPE1 `PP_PU_META_TYPE1_POS:`PP_PU_META_TID_POS+1
`define PP_PU_META_F_PAYLOAD_RANGE `PP_PU_META_F_PAYLOAD_NBITS-1:0
`define PP_PU_META_F_PAYLOAD_POS `PP_PU_META_F_PAYLOAD_NBITS+`PP_PU_META_TYPE1_POS
`define PP_PU_META_F_PAYLOAD `PP_PU_META_F_PAYLOAD_POS:`PP_PU_META_TYPE1_POS+1
`define PP_PU_META_T_PAYLOAD_RANGE `PP_PU_META_T_PAYLOAD_NBITS-1:0
`define PP_PU_META_T_PAYLOAD_POS `PP_PU_META_T_PAYLOAD_NBITS+`PP_PU_META_F_PAYLOAD_POS
`define PP_PU_META_T_PAYLOAD `PP_PU_META_T_PAYLOAD_POS:`PP_PU_META_F_PAYLOAD_POS+1

`define PU_QUEUE_PAYLOAD_LEN_NBITS `HOP_ID_NBITS
`define PU_QUEUE_PAYLOAD_PD_LEN_NBITS `PD_CHUNK_NBITS
`define PU_QUEUE_PAYLOAD_INST_LEN_NBITS `INST_CHUNK_NBITS
`define PU_QUEUE_PAYLOAD_BUF_PTR_NBITS `PIARB_BUF_PTR_NBITS
`define PU_QUEUE_PAYLOAD_INST_BUF_PTR_NBITS `PIARB_INST_BUF_PTR_NBITS
`define PU_QUEUE_PAYLOAD_PP_META_NBITS `PP_PIARB_META_NBITS
`define PU_QUEUE_PAYLOAD_NBITS `PU_QUEUE_PAYLOAD_PP_META_NBITS+`PU_QUEUE_PAYLOAD_INST_BUF_PTR_NBITS+`PU_QUEUE_PAYLOAD_BUF_PTR_NBITS+`PU_QUEUE_PAYLOAD_INST_LEN_NBITS+`PU_QUEUE_PAYLOAD_PD_LEN_NBITS+`PU_QUEUE_PAYLOAD_LEN_NBITS
`define PU_QUEUE_PAYLOAD_RANGE `PU_QUEUE_PAYLOAD_NBITS-1:0
`define PU_QUEUE_PAYLOAD_LEN_RANGE `PU_QUEUE_PAYLOAD_LEN_NBITS-1:0
`define PU_QUEUE_PAYLOAD_LEN_POS `PU_QUEUE_PAYLOAD_LEN_NBITS-1
`define PU_QUEUE_PAYLOAD_LEN `PU_QUEUE_PAYLOAD_LEN_POS:0
`define PU_QUEUE_PAYLOAD_PD_LEN_RANGE `PU_QUEUE_PAYLOAD_PD_LEN_NBITS-1:0
`define PU_QUEUE_PAYLOAD_PD_LEN_POS `PU_QUEUE_PAYLOAD_PD_LEN_NBITS+`PU_QUEUE_PAYLOAD_LEN_POS
`define PU_QUEUE_PAYLOAD_PD_LEN `PU_QUEUE_PAYLOAD_PD_LEN_POS:`PU_QUEUE_PAYLOAD_LEN_POS+1
`define PU_QUEUE_PAYLOAD_INST_LEN_RANGE `PU_QUEUE_PAYLOAD_INST_LEN_NBITS-1:0
`define PU_QUEUE_PAYLOAD_INST_LEN_POS `PU_QUEUE_PAYLOAD_INST_LEN_NBITS+`PU_QUEUE_PAYLOAD_PD_LEN_POS
`define PU_QUEUE_PAYLOAD_INST_LEN `PU_QUEUE_PAYLOAD_INST_LEN_POS:`PU_QUEUE_PAYLOAD_PD_LEN_POS+1
`define PU_QUEUE_PAYLOAD_BUF_PTR_RANGE `PU_QUEUE_PAYLOAD_BUF_PTR_NBITS-1:0
`define PU_QUEUE_PAYLOAD_BUF_PTR_POS `PU_QUEUE_PAYLOAD_BUF_PTR_NBITS+`PU_QUEUE_PAYLOAD_INST_LEN_POS
`define PU_QUEUE_PAYLOAD_BUF_PTR `PU_QUEUE_PAYLOAD_BUF_PTR_POS:`PU_QUEUE_PAYLOAD_INST_LEN_POS+1
`define PU_QUEUE_PAYLOAD_INST_BUF_PTR_RANGE `PU_QUEUE_PAYLOAD_INST_BUF_PTR_NBITS-1:0
`define PU_QUEUE_PAYLOAD_INST_BUF_PTR_POS `PU_QUEUE_PAYLOAD_INST_BUF_PTR_NBITS+`PU_QUEUE_PAYLOAD_BUF_PTR_POS
`define PU_QUEUE_PAYLOAD_INST_BUF_PTR `PU_QUEUE_PAYLOAD_INST_BUF_PTR_POS:`PU_QUEUE_PAYLOAD_BUF_PTR_POS+1
`define PU_QUEUE_PAYLOAD_PP_META_RANGE `PU_QUEUE_PAYLOAD_PP_META_NBITS-1:0
`define PU_QUEUE_PAYLOAD_PP_META_POS `PU_QUEUE_PAYLOAD_PP_META_NBITS+`PU_QUEUE_PAYLOAD_BUF_PTR_POS
`define PU_QUEUE_PAYLOAD_PP_META `PU_QUEUE_PAYLOAD_PP_META_POS:`PU_QUEUE_PAYLOAD_BUF_PTR_POS+1

`define PKT_DESC_DEPTH_NBITS 12
`define PKT_DESC_DEPTH (1<<`PKT_DESC_DEPTH_NBITS)

`define SCH_PKT_DESC_SRC_PORT_NBITS `PORT_ID_NBITS
`define SCH_PKT_DESC_DST_PORT_NBITS `PORT_ID_NBITS
`define SCH_PKT_DESC_PKT_LEN_NBITS `PACKET_LENGTH_NBITS
`define SCH_PKT_DESC_IDX_NBITS `PKT_DESC_DEPTH_NBITS
`define SCH_PKT_DESC_NBITS `SCH_PKT_DESC_IDX_NBITS+`SCH_PKT_DESC_PKT_LEN_NBITS+`SCH_PKT_DESC_DST_PORT_NBITS+`SCH_PKT_DESC_SRC_PORT_NBITS
`define SCH_PKT_DESC_RANGE `SCH_PKT_DESC_NBITS-1:0
`define SCH_PKT_DESC_SRC_PORT_RANGE `SCH_PKT_DESC_SRC_PORT_NBITS-1:0
`define SCH_PKT_DESC_SRC_PORT_POS `SCH_PKT_DESC_SRC_PORT_NBITS-1
`define SCH_PKT_DESC_SRC_PORT `SCH_PKT_DESC_SRC_PORT_POS:0
`define SCH_PKT_DESC_DST_PORT_RANGE `SCH_PKT_DESC_DST_PORT_NBITS-1:0
`define SCH_PKT_DESC_DST_PORT_POS `SCH_PKT_DESC_DST_PORT_NBITS+`SCH_PKT_DESC_SRC_PORT_POS
`define SCH_PKT_DESC_DST_PORT `SCH_PKT_DESC_DST_PORT_POS:`SCH_PKT_DESC_SRC_PORT_POS+1
`define SCH_PKT_DESC_PKT_LEN_RANGE `SCH_PKT_DESC_PKT_LEN_NBITS-1:0
`define SCH_PKT_DESC_PKT_LEN_POS `SCH_PKT_DESC_PKT_LEN_NBITS+`SCH_PKT_DESC_DST_PORT_POS
`define SCH_PKT_DESC_PKT_LEN `SCH_PKT_DESC_PKT_LEN_POS:`SCH_PKT_DESC_DST_PORT_POS+1
`define SCH_PKT_DESC_IDX_RANGE `SCH_PKT_DESC_IDX_NBITS-1:0
`define SCH_PKT_DESC_IDX_POS `SCH_PKT_DESC_IDX_NBITS+`SCH_PKT_DESC_PKT_LEN_POS
`define SCH_PKT_DESC_IDX `SCH_PKT_DESC_IDX_POS:`SCH_PKT_DESC_PKT_LEN_POS+1

`define PKT_DESC_QUEUE_NBITS `FIRST_LVL_QUEUE_ID_NBITS
`define PKT_DESC_CONN_NBITS `SECOND_LVL_QUEUE_ID_NBITS
`define PKT_DESC_CONN_GROUP_NBITS `THIRD_LVL_QUEUE_ID_NBITS
`define PKT_DESC_PORT_QUEUE_NBITS `FOURTH_LVL_QUEUE_ID_NBITS
`define PKT_DESC_SCH_DESC_NBITS `SCH_PKT_DESC_NBITS
`define PKT_DESC_NBITS `PKT_DESC_CONN_GROUP_NBITS+`PKT_DESC_CONN_NBITS+`PKT_DESC_QUEUE_NBITS+`PKT_DESC_PORT_QUEUE_NBITS+`PKT_DESC_SCH_DESC_NBITS
`define PKT_DESC_RANGE `PKT_DESC_NBITS-1:0
`define PKT_DESC_QUEUE_RANGE `PKT_DESC_QUEUE_NBITS-1:0
`define PKT_DESC_QUEUE_POS `PKT_DESC_QUEUE_NBITS-1
`define PKT_DESC_QUEUE `PKT_DESC_QUEUE_POS:0
`define PKT_DESC_CONN_RANGE `PKT_DESC_CONN_NBITS-1:0
`define PKT_DESC_CONN_POS `PKT_DESC_CONN_NBITS+`PKT_DESC_QUEUE_POS
`define PKT_DESC_CONN `PKT_DESC_CONN_POS:`PKT_DESC_QUEUE_POS+1
`define PKT_DESC_CONN_GROUP_RANGE `PKT_DESC_CONN_GROUP_NBITS-1:0
`define PKT_DESC_CONN_GROUP_POS `PKT_DESC_CONN_GROUP_NBITS+`PKT_DESC_CONN_POS
`define PKT_DESC_CONN_GROUP `PKT_DESC_CONN_GROUP_POS:`PKT_DESC_CONN_POS+1
`define PKT_DESC_PORT_QUEUE_RANGE `PKT_DESC_PORT_QUEUE_NBITS-1:0
`define PKT_DESC_PORT_QUEUE_POS `PKT_DESC_PORT_QUEUE_NBITS+`PKT_DESC_CONN_GROUP_POS
`define PKT_DESC_PORT_QUEUE `PKT_DESC_PORT_QUEUE_POS:`PKT_DESC_CONN_GROUP_POS+1
`define PKT_DESC_SCH_DESC_RANGE `PKT_DESC_SCH_DESC_NBITS-1:0
`define PKT_DESC_SCH_DESC_POS `PKT_DESC_SCH_DESC_NBITS+`PKT_DESC_PORT_QUEUE_POS
`define PKT_DESC_SCH_DESC `PKT_DESC_SCH_DESC_POS:`PKT_DESC_PORT_QUEUE_POS+1

`define ENQ_PKT_DESC_SRC_PORT_NBITS `PORT_ID_NBITS
`define ENQ_PKT_DESC_DST_PORT_NBITS `PORT_ID_NBITS
`define ENQ_PKT_DESC_BUF_PTR_NBITS `BUF_PTR_NBITS
`define ENQ_PKT_DESC_ED_CMD_NBITS `ENQ_ED_CMD_NBITS
`define ENQ_PKT_DESC_NBITS `ENQ_PKT_DESC_ED_CMD_NBITS+`ENQ_PKT_DESC_BUF_PTR_NBITS+`ENQ_PKT_DESC_DST_PORT_NBITS+`ENQ_PKT_DESC_SRC_PORT_NBITS
`define ENQ_PKT_DESC_RANGE `ENQ_PKT_DESC_NBITS-1:0
`define ENQ_PKT_DESC_SRC_PORT_RANGE `ENQ_PKT_DESC_SRC_PORT_NBITS-1:0
`define ENQ_PKT_DESC_SRC_PORT_POS `ENQ_PKT_DESC_SRC_PORT_NBITS-1
`define ENQ_PKT_DESC_SRC_PORT `ENQ_PKT_DESC_SRC_PORT_POS:0
`define ENQ_PKT_DESC_DST_PORT_RANGE `ENQ_PKT_DESC_DST_PORT_NBITS-1:0
`define ENQ_PKT_DESC_DST_PORT_POS `ENQ_PKT_DESC_DST_PORT_NBITS+`ENQ_PKT_DESC_SRC_PORT_POS
`define ENQ_PKT_DESC_DST_PORT `ENQ_PKT_DESC_DST_PORT_POS:`ENQ_PKT_DESC_SRC_PORT_POS+1
`define ENQ_PKT_DESC_BUF_PTR_RANGE `ENQ_PKT_DESC_BUF_PTR_NBITS-1:0
`define ENQ_PKT_DESC_BUF_PTR_POS `ENQ_PKT_DESC_BUF_PTR_NBITS+`ENQ_PKT_DESC_DST_PORT_POS
`define ENQ_PKT_DESC_BUF_PTR `ENQ_PKT_DESC_BUF_PTR_POS:`ENQ_PKT_DESC_DST_PORT_POS+1
`define ENQ_PKT_DESC_ED_CMD_RANGE `ENQ_PKT_DESC_ED_CMD_NBITS-1:0
`define ENQ_PKT_DESC_ED_CMD_POS `ENQ_PKT_DESC_ED_CMD_NBITS+`ENQ_PKT_DESC_BUF_PTR_POS
`define ENQ_PKT_DESC_ED_CMD `ENQ_PKT_DESC_ED_CMD_POS:`ENQ_PKT_DESC_BUF_PTR_POS+1

`define ASA_PROC_META_ED_CMD_NBITS `ENQ_ED_CMD_NBITS
`define ASA_PROC_META_BUF_PTR_NBITS `BUF_PTR_NBITS
`define ASA_PROC_META_FID_NBITS `FID_NBITS
`define ASA_PROC_META_TID_NBITS `TID_NBITS
`define ASA_PROC_META_TYPE1_NBITS 1
`define ASA_PROC_META_SRC_PORT_NBITS `PORT_ID_NBITS
`define ASA_PROC_META_DST_PORT_NBITS `PORT_ID_NBITS
`define ASA_PROC_META_IN_RCI_NBITS `RCI_NBITS
`define ASA_PROC_META_DOMAIN_ID_NBITS `DOMAIN_ID_NBITS
`define ASA_PROC_META_TIME_NBITS `PIARB_ASA_META_TIME_NBITS
`define ASA_PROC_META_DISCARD_NBITS 1
`define ASA_PROC_META_NBITS `ASA_PROC_META_DISCARD_NBITS+`ASA_PROC_META_TIME_NBITS+`ASA_PROC_META_DOMAIN_ID_NBITS+`ASA_PROC_META_IN_RCI_NBITS+`ASA_PROC_META_DST_PORT_NBITS+`ASA_PROC_META_SRC_PORT_NBITS+`ASA_PROC_META_TYPE1_NBITS+`ASA_PROC_META_TID_NBITS+`ASA_PROC_META_FID_NBITS+`ASA_PROC_META_BUF_PTR_NBITS+`ASA_PROC_META_ED_CMD_NBITS
`define ASA_PROC_META_RANGE `ASA_PROC_META_NBITS-1:0
`define ASA_PROC_META_ED_CMD_RANGE `ASA_PROC_META_ED_CMD_NBITS-1:0
`define ASA_PROC_META_ED_CMD_POS `ASA_PROC_META_ED_CMD_NBITS-1
`define ASA_PROC_META_ED_CMD `ASA_PROC_META_ED_CMD_POS:0
`define ASA_PROC_META_BUF_PTR_RANGE `ASA_PROC_META_BUF_PTR_NBITS-1:0
`define ASA_PROC_META_BUF_PTR_POS `ASA_PROC_META_BUF_PTR_NBITS+`ASA_PROC_META_ED_CMD_POS
`define ASA_PROC_META_BUF_PTR `ASA_PROC_META_BUF_PTR_POS:`ASA_PROC_META_ED_CMD_POS+1
`define ASA_PROC_META_FID_RANGE `ASA_PROC_META_FID_NBITS-1:0
`define ASA_PROC_META_FID_POS `ASA_PROC_META_FID_NBITS+`ASA_PROC_META_BUF_PTR_POS
`define ASA_PROC_META_FID `ASA_PROC_META_FID_POS:`ASA_PROC_META_BUF_PTR_POS+1
`define ASA_PROC_META_TID_RANGE `ASA_PROC_META_TID_NBITS-1:0
`define ASA_PROC_META_TID_POS `ASA_PROC_META_TID_NBITS+`ASA_PROC_META_FID_POS
`define ASA_PROC_META_TID `ASA_PROC_META_TID_POS:`ASA_PROC_META_FID_POS+1
`define ASA_PROC_META_TYPE1_RANGE `ASA_PROC_META_TYPE1_NBITS-1:0
`define ASA_PROC_META_TYPE1_POS `ASA_PROC_META_TYPE1_NBITS+`ASA_PROC_META_TID_POS
`define ASA_PROC_META_TYPE1 `ASA_PROC_META_TYPE1_POS:`ASA_PROC_META_TID_POS+1
`define ASA_PROC_META_SRC_PORT_RANGE `ASA_PROC_META_SRC_PORT_NBITS-1:0
`define ASA_PROC_META_SRC_PORT_POS `ASA_PROC_META_SRC_PORT_NBITS+`ASA_PROC_META_TYPE1_POS
`define ASA_PROC_META_SRC_PORT `ASA_PROC_META_SRC_PORT_POS:`ASA_PROC_META_TYPE1_POS+1
`define ASA_PROC_META_DST_PORT_RANGE `ASA_PROC_META_DST_PORT_NBITS-1:0
`define ASA_PROC_META_DST_PORT_POS `ASA_PROC_META_DST_PORT_NBITS+`ASA_PROC_META_SRC_PORT_POS
`define ASA_PROC_META_DST_PORT `ASA_PROC_META_DST_PORT_POS:`ASA_PROC_META_SRC_PORT_POS+1
`define ASA_PROC_META_IN_RCI_RANGE `ASA_PROC_META_IN_RCI_NBITS-1:0
`define ASA_PROC_META_IN_RCI_POS `ASA_PROC_META_IN_RCI_NBITS+`ASA_PROC_META_DST_PORT_POS
`define ASA_PROC_META_IN_RCI `ASA_PROC_META_IN_RCI_POS:`ASA_PROC_META_DST_PORT_POS+1
`define ASA_PROC_META_DOMAIN_ID_RANGE `ASA_PROC_META_DOMAIN_ID_NBITS-1:0
`define ASA_PROC_META_DOMAIN_ID_POS `ASA_PROC_META_DOMAIN_ID_NBITS+`ASA_PROC_META_IN_RCI_POS
`define ASA_PROC_META_DOMAIN_ID `ASA_PROC_META_DOMAIN_ID_POS:`ASA_PROC_META_IN_RCI_POS+1
`define ASA_PROC_META_TIME_RANGE `ASA_PROC_META_TIME_NBITS-1:0
`define ASA_PROC_META_TIME_POS `ASA_PROC_META_TIME_NBITS+`ASA_PROC_META_DOMAIN_ID_POS
`define ASA_PROC_META_TIME `ASA_PROC_META_TIME_POS:`ASA_PROC_META_DOMAIN_ID_POS+1
`define ASA_PROC_META_DISCARD_RANGE `ASA_PROC_META_DISCARD_NBITS-1:0
`define ASA_PROC_META_DISCARD_POS `ASA_PROC_META_DISCARD_NBITS+`ASA_PROC_META_TIME_POS
`define ASA_PROC_META_DISCARD `ASA_PROC_META_DISCARD_POS:`ASA_PROC_META_TIME_POS+1

`define RAS_FLAG_UPPD_NBITS 1
`define RAS_FLAG_UPPP_NBITS 1
`define RAS_FLAG_UFDAST_NBITS 3
`define RAS_FLAG_EAST_NBITS 3
`define RAS_FLAG_NFASCF_NBITS 2
`define RAS_FLAG_PTR_NBITS 16
`define RAS_FLAG_NBITS `RAS_FLAG_EAST_NBITS+`RAS_FLAG_UFDAST_NBITS+`RAS_FLAG_UPPP_NBITS+`RAS_FLAG_UPPD_NBITS+`RAS_FLAG_NFASCF_NBITS+`RAS_FLAG_PTR_NBITS
`define RAS_FLAG_RANGE `RAS_FLAG_NBITS-1:0
`define RAS_FLAG_UPPD_RANGE `RAS_FLAG_UPPD_NBITS-1:0
`define RAS_FLAG_UPPD_POS `RAS_FLAG_UPPD_NBITS-1
`define RAS_FLAG_UPPD `RAS_FLAG_UPPD_POS:0
`define RAS_FLAG_UPPP_RANGE `RAS_FLAG_UPPP_NBITS-1:0
`define RAS_FLAG_UPPP_POS `RAS_FLAG_UPPP_NBITS+`RAS_FLAG_UPPD_POS
`define RAS_FLAG_UPPP `RAS_FLAG_UPPP_POS:`RAS_FLAG_UPPD_POS+1
`define RAS_FLAG_UFDAST_RANGE `RAS_FLAG_UFDAST_NBITS-1:0
`define RAS_FLAG_UFDAST_POS `RAS_FLAG_UFDAST_NBITS+`RAS_FLAG_UPPP_POS
`define RAS_FLAG_UFDAST `RAS_FLAG_UFDAST_POS:`RAS_FLAG_UPPP_POS+1
`define RAS_FLAG_EAST_RANGE `RAS_FLAG_EAST_NBITS-1:0
`define RAS_FLAG_EAST_POS `RAS_FLAG_EAST_NBITS+`RAS_FLAG_UFDAST_POS
`define RAS_FLAG_EAST `RAS_FLAG_EAST_POS:`RAS_FLAG_UFDAST_POS+1
`define RAS_FLAG_NFASCF_RANGE `RAS_FLAG_NFASCF_NBITS-1:0
`define RAS_FLAG_NFASCF_POS `RAS_FLAG_NFASCF_NBITS+`RAS_FLAG_EAST_POS
`define RAS_FLAG_NFASCF `RAS_FLAG_NFASCF_POS:`RAS_FLAG_EAST_POS+1
`define RAS_FLAG_PTR_RANGE `RAS_FLAG_PTR_NBITS-1:0
`define RAS_FLAG_PTR_POS `RAS_FLAG_PTR_NBITS+`RAS_FLAG_NFASCF_POS
`define RAS_FLAG_PTR `RAS_FLAG_PTR_POS:`RAS_FLAG_NFASCF_POS+1

`define RAS_NBITS (`RAS_FLAG_NBITS+(1+`SCI_NBITS)*9)

`define DECR_BLOCK_ADDR_LSB             20 
`define DECR_BLOCK_ADDR             12'd0
`define DECR_MEM_ADDR_MSB             `DECR_BLOCK_ADDR_LSB-1 
`define DECR_MEM_ADDR_LSB             `RCI_VALUE_DEPTH_NBITS+6
`define DECR_MEM_ADDR_RANGE             `DECR_MEM_ADDR_MSB:`DECR_MEM_ADDR_LSB 

`define ENCR_BLOCK_ADDR_LSB             20 
`define ENCR_BLOCK_ADDR             12'd1
`define ENCR_MEM_ADDR_MSB             `ENCR_BLOCK_ADDR_LSB-1 
`define ENCR_MEM_ADDR_LSB             `EEKEY_VALUE_DEPTH_NBITS+6
`define ENCR_MEM_ADDR_RANGE             `ENCR_MEM_ADDR_MSB:`ENCR_MEM_ADDR_LSB 

`define TM_BLOCK_ADDR_LSB             20 
`define TM_BLOCK_ADDR             12'd2
`define TM_MEM_ADDR_MSB             `TM_BLOCK_ADDR_LSB-1 
`define TM_MEM_ADDR_LSB             `FIRST_LVL_QUEUE_ID_NBITS+2
`define TM_MEM_ADDR_RANGE             `TM_MEM_ADDR_MSB:`TM_MEM_ADDR_LSB 

`define ASA_BLOCK_ADDR_LSB             20 
`define ASA_BLOCK_ADDR             12'd3
`define ASA_MEM_ADDR_MSB             `ASA_BLOCK_ADDR_LSB-1 
`define ASA_MEM_ADDR_LSB             `RCI_NBITS+2
`define ASA_MEM_ADDR_RANGE             `ASA_MEM_ADDR_MSB:`ASA_MEM_ADDR_LSB 

`define CLASSIFIER_BLOCK_ADDR_LSB             20 
`define CLASSIFIER_BLOCK_ADDR             12'd4
`define CLASSIFIER_MEM_ADDR_MSB             `CLASSIFIER_BLOCK_ADDR_LSB-1 
`define CLASSIFIER_MEM_ADDR_LSB             `FLOW_HASH_TABLE_DEPTH_NBITS+4
`define CLASSIFIER_MEM_ADDR_RANGE             `CLASSIFIER_MEM_ADDR_MSB:`CLASSIFIER_MEM_ADDR_LSB 

`define IRL_BLOCK_ADDR_LSB             20 
`define IRL_BLOCK_ADDR             12'd5
`define IRL_MEM_ADDR_MSB             `IRL_BLOCK_ADDR_LSB-1 
`define IRL_MEM_ADDR_LSB             `LIMITER_NBITS+2
`define IRL_MEM_ADDR_RANGE             `IRL_MEM_ADDR_MSB:`IRL_MEM_ADDR_LSB 

`define PIARB_BLOCK_ADDR_LSB             20 
`define PIARB_BLOCK_ADDR             12'd6
`define PIARB_MEM_ADDR_MSB             `PIARB_BLOCK_ADDR_LSB-1 
`define PIARB_MEM_ADDR_LSB             `TID_NBITS+2
`define PIARB_MEM_ADDR_RANGE             `PIARB_MEM_ADDR_MSB:`PIARB_MEM_ADDR_LSB 

`define PU_BLOCK_ADDR_LSB             20 
`define PU_BLOCK_ADDR             12'd7
`define PU_MEM_ADDR_MSB             `PU_BLOCK_ADDR_LSB-1 
`define PU_MEM_ADDR_LSB             `SCI_NBITS+`CONNECTION_CONTEXT_DEPTH_NBITS+2
`define PU_MEM_ADDR_RANGE             `PU_MEM_ADDR_MSB:`PU_MEM_ADDR_LSB 

`define REG_BLOCK_ADDR 12'd8

`define ECDSA_BLOCK_ADDR_LSB             20 
`define BM_BLOCK_ADDR_LSB             20 
`define BM_BLOCK_ADDR             12'd9

`define BM_REG_BLOCK_ADDR_LSB             8 
`define BM_REG_BLOCK_ADDR             {`REG_BLOCK_ADDR, {(`BM_BLOCK_ADDR_LSB-`BM_REG_BLOCK_ADDR_LSB-9){1'b0}}, 9'd0}
`define BM_REG_ADDR_RANGE             `BM_BLOCK_ADDR_LSB-1:`PIO_ADDR_LSB 

`define ENCR_REG_BLOCK_ADDR_LSB             8 
`define ENCR_REG_BLOCK_ADDR             {`REG_BLOCK_ADDR, {(`ENCR_BLOCK_ADDR_LSB-`ENCR_REG_BLOCK_ADDR_LSB-9){1'b0}}, 9'd1}
`define ENCR_REG_ADDR_RANGE             `ENCR_REG_BLOCK_ADDR_LSB-1:`PIO_ADDR_LSB 

`define ASA_REG_BLOCK_ADDR_LSB             8 
`define ASA_REG_BLOCK_ADDR             {`REG_BLOCK_ADDR, {(`ASA_BLOCK_ADDR_LSB-`ASA_REG_BLOCK_ADDR_LSB-9){1'b0}}, 9'd2}
`define ASA_REG_ADDR_RANGE             `ASA_REG_BLOCK_ADDR_LSB-1:`PIO_ADDR_LSB 

`define CLASSIFIER_REG_BLOCK_ADDR_LSB             8 
`define CLASSIFIER_REG_BLOCK_ADDR             {`REG_BLOCK_ADDR, {(`CLASSIFIER_BLOCK_ADDR_LSB-`CLASSIFIER_REG_BLOCK_ADDR_LSB-9){1'b0}}, 9'd3}
`define CLASSIFIER_REG_ADDR_RANGE             `CLASSIFIER_REG_BLOCK_ADDR_LSB-1:`PIO_ADDR_LSB 

`define ECDSA_REG_BLOCK_ADDR_LSB             8 
`define ECDSA_REG_BLOCK_ADDR             {`REG_BLOCK_ADDR, {(`ECDSA_BLOCK_ADDR_LSB-`ECDSA_REG_BLOCK_ADDR_LSB-9){1'b0}}, 9'd4}
`define ECDSA_REG_ADDR_RANGE             `ECDSA_REG_BLOCK_ADDR_LSB-1:`PIO_ADDR_LSB 

`define BM_FREEB_INIT            6'd0 
`define BM_FREEB_RD_COUNT            6'd1 
`define BM_FREEB_WR_COUNT            6'd2 
`define BM_LL_RD_COUNT            6'd3 
`define BM_LL_WR_COUNT            6'd4 
`define BM_DT_ALPHA            6'd5 

`define ENCR_MAC_SA_LSB            6'd0 
`define ENCR_MAC_SA_MSB            6'd1 
`define ENCR_IPSEC_IV_LSB            6'd2 
`define ENCR_IPSEC_IV_MSB            6'd3 
`define ENCR_GRE_HEADER            6'd4 
`define ENCR_ID_TTL_DSCP            6'd5 
`define ENCR_FLOW_LABEL            6'd6 
`define ENCR_IN_MAC_SA_LSB            6'd7 
`define ENCR_IN_MAC_SA_MSB            6'd8 
`define ENCR_IN_MAC_DA_LSB            6'd9 
`define ENCR_IN_MAC_DA_MSB            6'd10 
`define ENCR_IN_VLAN            6'd11 

`define ASA_DEFAULT_SUB_EXP_TIME            6'd0 
`define ASA_SUPERVISOR_SCI            6'd1 
`define ASA_CLASS2PRI            6'd2 

`define CLASSIFIER_AGING_TIME            6'd0 

`define ECDSA_DEFAULT_EXP_TIME            6'd0 

`define TM_QUEUE_ASSOCIATION             6'd15
`define TM_QUEUE_PROFILE0             6'd8
`define TM_WDRR_QUANTUM0             6'd9
`define TM_SHAPING_PROFILE_CIR0             6'd10
`define TM_SHAPING_PROFILE_EIR0             6'd11
`define TM_WDRR_SCH_CTRL0             6'd12
`define TM_FILL_TB_DST0             6'd13
`define TM_PRI_SCH_CTRL00             6'd0
`define TM_PRI_SCH_CTRL01             6'd1
`define TM_PRI_SCH_CTRL02             6'd2
`define TM_PRI_SCH_CTRL03             6'd3
`define TM_PRI_SCH_CTRL04             6'd4
`define TM_PRI_SCH_CTRL05             6'd5
`define TM_PRI_SCH_CTRL06             6'd6
`define TM_PRI_SCH_CTRL07             6'd7
`define TM_QUEUE_PROFILE1             6'd24
`define TM_WDRR_QUANTUM1             6'd25
`define TM_SHAPING_PROFILE_CIR1             6'd26
`define TM_SHAPING_PROFILE_EIR1             6'd27
`define TM_WDRR_SCH_CTRL1             6'd28
`define TM_FILL_TB_DST1             6'd29
`define TM_PRI_SCH_CTRL10             6'd16
`define TM_PRI_SCH_CTRL11             6'd17
`define TM_PRI_SCH_CTRL12             6'd18
`define TM_PRI_SCH_CTRL13             6'd19
`define TM_PRI_SCH_CTRL14             6'd20
`define TM_PRI_SCH_CTRL15             6'd21
`define TM_PRI_SCH_CTRL16             6'd22
`define TM_PRI_SCH_CTRL17             6'd23
`define TM_QUEUE_PROFILE2             6'd40
`define TM_WDRR_QUANTUM2             6'd41
`define TM_SHAPING_PROFILE_CIR2             6'd42
`define TM_SHAPING_PROFILE_EIR2             6'd43
`define TM_WDRR_SCH_CTRL2             6'd44
`define TM_FILL_TB_DST2             6'd45
`define TM_PRI_SCH_CTRL20             6'd32
`define TM_PRI_SCH_CTRL21             6'd33
`define TM_PRI_SCH_CTRL22             6'd34
`define TM_PRI_SCH_CTRL23             6'd35
`define TM_PRI_SCH_CTRL24             6'd36
`define TM_PRI_SCH_CTRL25             6'd37
`define TM_PRI_SCH_CTRL26             6'd38
`define TM_PRI_SCH_CTRL27             6'd39
`define TM_QUEUE_PROFILE3             6'd56
`define TM_WDRR_QUANTUM3             6'd57
`define TM_SHAPING_PROFILE_CIR3             6'd58
`define TM_SHAPING_PROFILE_EIR3             6'd59
`define TM_WDRR_SCH_CTRL3             6'd60
`define TM_FILL_TB_DST3             6'd61
`define TM_PRI_SCH_CTRL30             6'd48
`define TM_PRI_SCH_CTRL31             6'd49
`define TM_PRI_SCH_CTRL32             6'd50
`define TM_PRI_SCH_CTRL33             6'd51
`define TM_PRI_SCH_CTRL34             6'd52
`define TM_PRI_SCH_CTRL35             6'd53
`define TM_PRI_SCH_CTRL36             6'd54
`define TM_PRI_SCH_CTRL37             6'd55

`define IRL_LIMITING_PROFILE_CIR           2'd0
`define IRL_LIMITING_PROFILE_EIR           2'd2
`define IRL_FILL_TB_SRC           2'd3

`define CLASSIFIER_FLOW_HASH_TABLE           2'd0
`define CLASSIFIER_TOPIC_HASH_TABLE           2'd2

`define DECR_RCI_HASH_TABLE           2'd0
`define DECR_RCI_VALUE           2'd1
`define DECR_EKEY_HASH_TABLE           2'd2
`define DECR_EKEY_VALUE           2'd3

`define ENCR_TUNNEL_HASH_TABLE           2'd0
`define ENCR_TUNNEL_VALUE           2'd1
`define ENCR_EEKEY_HASH_TABLE           2'd2
`define ENCR_EEKEY_VALUE           2'd3

`define ECDSA_TOPIC_POLICY 2'd0

`define PIARB_TOPIC_VALUE 2'd0

`define HASH(FUNC_NAME, KEY_NBITS, HASH_NBITS) \
function logic [HASH_NBITS-1:0] FUNC_NAME (input [KEY_NBITS-1:0] key);\
logic [(KEY_NBITS/HASH_NBITS)-1:0] key_div[HASH_NBITS-1:0]; 	\
logic [HASH_NBITS-1:0] pre_hash_value;	\
		\
integer i, j; \
begin \
		\
	for (i=0; i<HASH_NBITS; i++)	\
		for (j=0; j<(KEY_NBITS/HASH_NBITS); j++) \
			key_div[i][j] = key[j*HASH_NBITS+i];	\
			\
	for (i=0; i<HASH_NBITS; i++)	\
		pre_hash_value[i] = ^key_div[i];	\
		\
	FUNC_NAME = (KEY_NBITS%HASH_NBITS)==0?pre_hash_value:pre_hash_value^key[KEY_NBITS-1:KEY_NBITS-1-(KEY_NBITS%HASH_NBITS)-1];	\
end \
endfunction \

`define TRANSPOSE(FUNC_NAME, KEY_NBITS) \
function logic [KEY_NBITS-1:0] FUNC_NAME (input [KEY_NBITS-1:0] key);\
integer i; \
begin \
		\
	for (i=0; i<KEY_NBITS+1; i++)	\
		FUNC_NAME[i] = key[KEY_NBITS-1-i];	\
end \
endfunction \

`endif
