package core_test_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import special_packet_pkg::*;
  import mac_agent_pkg::*;
  import dma_agent_pkg::*;
  import pio_wr_agent_pkg::*;
  import pio_rd_agent_pkg::*;
  import core_env_pkg::*;

  `include "bay_test_base.svh"
  `include "core_test_base.svh"
  `include "core_test_first.svh"
  `include "core_test_second.svh"
  `include "core_test_third.svh"
  `include "core_test_fourth.svh"
  `include "core_test_fifth.svh"
  `include "core_test_sixth.svh"
  `include "core_test_seventh.svh"
  `include "core_test_pp0.svh"
  `include "core_test_pp1.svh"
  `include "core_test_pp2.svh"
  `include "core_test_pp3.svh"
  `include "core_test_pp4.svh"
  `include "core_test_pp5.svh"
  `include "core_test_pp6.svh"
  `include "core_test_pp7.svh"
  `include "core_test_pp8.svh"
  `include "core_test_pp9.svh"
  `include "core_test_pp10.svh"
  `include "core_test_pp11.svh"
  `include "core_test_pp12.svh"
  `include "core_test_pp13.svh"
  `include "core_test_pu0.svh"

endpackage
