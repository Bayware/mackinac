/* (c) 2017 Bayware, Inc.
//
//   Project: Mackinac
//   Module:  class_pkg.sv
//   Owner:   G Walter
//   Date:    10/27/17
//
//   Summary:  package for classifier block-level tb & design
*/

package class_pkg;
    typedef bit [ 31:0 ] uint32_t;
    typedef enum { FAIL, PASS } pf_e;

endpackage
