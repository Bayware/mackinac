package pio_rd_agent_pkg ;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "pio_rd_config.svh"
  `include "pio_rd_transaction.svh"
  `include "pio_rd_driver.svh"
  `include "pio_rd_monitor.svh"
  `include "pio_rd_agent.svh"
  `include "pio_rd_sequence.svh"

endpackage
