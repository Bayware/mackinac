package pio_wr_agent_pkg ;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import ral_pkg::*;

  `include "pio_wr_config.svh"
  `include "pio_wr_transaction.svh"
  `include "pio_wr_driver.svh"
  `include "pio_wr_monitor.svh"
  `include "pio_wr_adapter.svh"
  `include "pio_wr_agent.svh"
  `include "pio_wr_sequence.svh"
  `include "pio_wr_sequence_ral.svh"

endpackage
